module mux_2_1_27_bits (out, in_0, in_1, select);
output	[26:0]	out ;
input	[26:0]	in_0, in_1 ;
input			select ;

bufif0		nb_00	(out[00], in_0[00], select) ;
bufif0		nb_01	(out[01], in_0[01], select) ;
bufif0		nb_02	(out[02], in_0[02], select) ;
bufif0		nb_03	(out[03], in_0[03], select) ;
bufif0		nb_04	(out[04], in_0[04], select) ;
bufif0		nb_05	(out[05], in_0[05], select) ;
bufif0		nb_06	(out[06], in_0[06], select) ;
bufif0		nb_07	(out[07], in_0[07], select) ;
bufif0		nb_08	(out[08], in_0[08], select) ;
bufif0		nb_09	(out[09], in_0[09], select) ;
bufif0		nb_10	(out[10], in_0[10], select) ;
bufif0		nb_11	(out[11], in_0[11], select) ;
bufif0		nb_12	(out[12], in_0[12], select) ;
bufif0		nb_13	(out[13], in_0[13], select) ;
bufif0		nb_14	(out[14], in_0[14], select) ;
bufif0		nb_15	(out[15], in_0[15], select) ;
bufif0		nb_16	(out[16], in_0[16], select) ;
bufif0		nb_17	(out[17], in_0[17], select) ;
bufif0		nb_18	(out[18], in_0[18], select) ;
bufif0		nb_19	(out[19], in_0[19], select) ;
bufif0		nb_20	(out[20], in_0[20], select) ;
bufif0		nb_21	(out[21], in_0[21], select) ;
bufif0		nb_22	(out[22], in_0[22], select) ;
bufif0		nb_23	(out[23], in_0[23], select) ;
bufif0		nb_24	(out[24], in_0[24], select) ;
bufif0		nb_25	(out[25], in_0[25], select) ;
bufif0		nb_26	(out[26], in_0[26], select) ;

bufif1		b_00	(out[00], in_1[00], select) ;
bufif1		b_01	(out[01], in_1[01], select) ;
bufif1		b_02	(out[02], in_1[02], select) ;
bufif1		b_03	(out[03], in_1[03], select) ;
bufif1		b_04	(out[04], in_1[04], select) ;
bufif1		b_05	(out[05], in_1[05], select) ;
bufif1		b_06	(out[06], in_1[06], select) ;
bufif1		b_07	(out[07], in_1[07], select) ;
bufif1		b_08	(out[08], in_1[08], select) ;
bufif1		b_09	(out[09], in_1[09], select) ;
bufif1		b_10	(out[10], in_1[10], select) ;
bufif1		b_11	(out[11], in_1[11], select) ;
bufif1		b_12	(out[12], in_1[12], select) ;
bufif1		b_13	(out[13], in_1[13], select) ;
bufif1		b_14	(out[14], in_1[14], select) ;
bufif1		b_15	(out[15], in_1[15], select) ;
bufif1		b_16	(out[16], in_1[16], select) ;
bufif1		b_17	(out[17], in_1[17], select) ;
bufif1		b_18	(out[18], in_1[18], select) ;
bufif1		b_19	(out[19], in_1[19], select) ;
bufif1		b_20	(out[20], in_1[20], select) ;
bufif1		b_21	(out[21], in_1[21], select) ;
bufif1		b_22	(out[22], in_1[22], select) ;
bufif1		b_23	(out[23], in_1[23], select) ;
bufif1		b_24	(out[24], in_1[24], select) ;
bufif1		b_25	(out[25], in_1[25], select) ;
bufif1		b_26	(out[26], in_1[26], select) ;

endmodule // mux_2_1
