module ShiftRight24(X,shamt,Y);
input [7:0] shamt;
input [23:0] X;
output wire [23:0] Y;
wire  [24:0] en;

Decoder24 D0(shamt,en);
bufif1 (Y[0],X[0],en[0]);
bufif1 (Y[0],X[1],en[1]);
bufif1 (Y[0],X[2],en[2]);
bufif1 (Y[0],X[3],en[3]); 
bufif1 (Y[0],X[4],en[4]);
bufif1 (Y[0],X[5],en[5]);
bufif1 (Y[0],X[6],en[6]);
bufif1 (Y[0],X[7],en[7]);
bufif1 (Y[0],X[8],en[8]);
bufif1 (Y[0],X[9],en[9]);
bufif1 (Y[0],X[10],en[10]);
bufif1 (Y[0],X[11],en[11]);
bufif1 (Y[0],X[12],en[12]);
bufif1 (Y[0],X[13],en[13]);
bufif1 (Y[0],X[14],en[14]);
bufif1 (Y[0],X[15],en[15]);
bufif1 (Y[0],X[16],en[16]);
bufif1 (Y[0],X[17],en[17]);
bufif1 (Y[0],X[18],en[18]);
bufif1 (Y[0],X[19],en[19]);
bufif1 (Y[0],X[20],en[20]);
bufif1 (Y[0],X[21],en[21]);
bufif1 (Y[0],X[22],en[22]);
bufif1 (Y[0],X[23],en[23]);

bufif1 (Y[1],X[1],en[0]);
bufif1 (Y[1],X[2],en[1]);
bufif1 (Y[1],X[3],en[2]);
bufif1 (Y[1],X[4],en[3]);
bufif1 (Y[1],X[5],en[4]);
bufif1 (Y[1],X[6],en[5]);
bufif1 (Y[1],X[7],en[6]);
bufif1 (Y[1],X[8],en[7]);
bufif1 (Y[1],X[9],en[8]);
bufif1 (Y[1],X[10],en[9]);
bufif1 (Y[1],X[11],en[10]);
bufif1 (Y[1],X[12],en[11]);
bufif1 (Y[1],X[13],en[12]);
bufif1 (Y[1],X[14],en[13]);
bufif1 (Y[1],X[15],en[14]);
bufif1 (Y[1],X[16],en[15]);
bufif1 (Y[1],X[17],en[16]);
bufif1 (Y[1],X[18],en[17]);
bufif1 (Y[1],X[19],en[18]);
bufif1 (Y[1],X[20],en[19]);
bufif1 (Y[1],X[21],en[20]);
bufif1 (Y[1],X[22],en[21]);
bufif1 (Y[1],X[23],en[22]);

bufif1 (Y[2],X[2],en[0]);
bufif1 (Y[2],X[3],en[1]);
bufif1 (Y[2],X[4],en[2]);
bufif1 (Y[2],X[5],en[3]);
bufif1 (Y[2],X[6],en[4]);
bufif1 (Y[2],X[7],en[5]);
bufif1 (Y[2],X[8],en[6]);
bufif1 (Y[2],X[9],en[7]);
bufif1 (Y[2],X[10],en[8]);
bufif1 (Y[2],X[11],en[9]);
bufif1 (Y[2],X[12],en[10]);
bufif1 (Y[2],X[13],en[11]);
bufif1 (Y[2],X[14],en[12]);
bufif1 (Y[2],X[15],en[13]);
bufif1 (Y[2],X[16],en[14]);
bufif1 (Y[2],X[17],en[15]);
bufif1 (Y[2],X[18],en[16]);
bufif1 (Y[2],X[19],en[17]);
bufif1 (Y[2],X[20],en[18]);
bufif1 (Y[2],X[21],en[19]);
bufif1 (Y[2],X[22],en[20]);
bufif1 (Y[2],X[23],en[21]);

bufif1 (Y[3],X[3],en[0]);
bufif1 (Y[3],X[4],en[1]);
bufif1 (Y[3],X[5],en[2]);
bufif1 (Y[3],X[6],en[3]);
bufif1 (Y[3],X[7],en[4]);
bufif1 (Y[3],X[8],en[5]);
bufif1 (Y[3],X[9],en[6]);
bufif1 (Y[3],X[10],en[7]);
bufif1 (Y[3],X[11],en[8]);
bufif1 (Y[3],X[12],en[9]);
bufif1 (Y[3],X[13],en[10]);
bufif1 (Y[3],X[14],en[11]);
bufif1 (Y[3],X[15],en[12]);
bufif1 (Y[3],X[16],en[13]);
bufif1 (Y[3],X[17],en[14]);
bufif1 (Y[3],X[18],en[15]);
bufif1 (Y[3],X[19],en[16]);
bufif1 (Y[3],X[20],en[17]);
bufif1 (Y[3],X[21],en[18]);
bufif1 (Y[3],X[22],en[19]);
bufif1 (Y[3],X[23],en[20]);

bufif1 (Y[4],X[4],en[0]);
bufif1 (Y[4],X[5],en[1]);
bufif1 (Y[4],X[6],en[2]);
bufif1 (Y[4],X[7],en[3]);
bufif1 (Y[4],X[8],en[4]);
bufif1 (Y[4],X[9],en[5]);
bufif1 (Y[4],X[10],en[6]);
bufif1 (Y[4],X[11],en[7]);
bufif1 (Y[4],X[12],en[8]);
bufif1 (Y[4],X[13],en[9]);
bufif1 (Y[4],X[14],en[10]);
bufif1 (Y[4],X[15],en[11]);
bufif1 (Y[4],X[16],en[12]);
bufif1 (Y[4],X[17],en[13]);
bufif1 (Y[4],X[18],en[14]);
bufif1 (Y[4],X[19],en[15]);
bufif1 (Y[4],X[20],en[16]);
bufif1 (Y[4],X[21],en[17]);
bufif1 (Y[4],X[22],en[18]);
bufif1 (Y[4],X[23],en[19]);

bufif1 (Y[5],X[5],en[0]);
bufif1 (Y[5],X[6],en[1]);
bufif1 (Y[5],X[7],en[2]);
bufif1 (Y[5],X[8],en[3]);
bufif1 (Y[5],X[9],en[4]);
bufif1 (Y[5],X[10],en[5]);
bufif1 (Y[5],X[11],en[6]);
bufif1 (Y[5],X[12],en[7]);
bufif1 (Y[5],X[13],en[8]);
bufif1 (Y[5],X[14],en[9]);
bufif1 (Y[5],X[15],en[10]);
bufif1 (Y[5],X[16],en[11]);
bufif1 (Y[5],X[17],en[12]);
bufif1 (Y[5],X[18],en[13]);
bufif1 (Y[5],X[19],en[14]);
bufif1 (Y[5],X[20],en[15]);
bufif1 (Y[5],X[21],en[16]);
bufif1 (Y[5],X[22],en[17]);
bufif1 (Y[5],X[23],en[18]);


bufif1 (Y[6],X[6],en[0]);
bufif1 (Y[6],X[7],en[1]);
bufif1 (Y[6],X[8],en[2]);
bufif1 (Y[6],X[9],en[3]);
bufif1 (Y[6],X[10],en[4]);
bufif1 (Y[6],X[11],en[5]);
bufif1 (Y[6],X[12],en[6]);
bufif1 (Y[6],X[13],en[7]);
bufif1 (Y[6],X[14],en[8]);
bufif1 (Y[6],X[15],en[9]);
bufif1 (Y[6],X[16],en[10]);
bufif1 (Y[6],X[17],en[11]);
bufif1 (Y[6],X[18],en[12]);
bufif1 (Y[6],X[19],en[13]);
bufif1 (Y[6],X[20],en[14]);
bufif1 (Y[6],X[21],en[15]);
bufif1 (Y[6],X[22],en[16]);
bufif1 (Y[6],X[23],en[17]);

bufif1 (Y[7],X[7],en[0]);
bufif1 (Y[7],X[8],en[1]);
bufif1 (Y[7],X[9],en[2]);
bufif1 (Y[7],X[10],en[3]);
bufif1 (Y[7],X[11],en[4]);
bufif1 (Y[7],X[12],en[5]);
bufif1 (Y[7],X[13],en[6]);
bufif1 (Y[7],X[14],en[7]);
bufif1 (Y[7],X[15],en[8]);
bufif1 (Y[7],X[16],en[9]);
bufif1 (Y[7],X[17],en[10]);
bufif1 (Y[7],X[18],en[11]);
bufif1 (Y[7],X[19],en[12]);
bufif1 (Y[7],X[20],en[13]);
bufif1 (Y[7],X[21],en[14]);
bufif1 (Y[7],X[22],en[15]);
bufif1 (Y[7],X[23],en[16]);

bufif1 (Y[8],X[8],en[0]);
bufif1 (Y[8],X[9],en[1]);
bufif1 (Y[8],X[10],en[2]);
bufif1 (Y[8],X[11],en[3]);
bufif1 (Y[8],X[12],en[4]);
bufif1 (Y[8],X[13],en[5]);
bufif1 (Y[8],X[14],en[6]);
bufif1 (Y[8],X[15],en[7]);
bufif1 (Y[8],X[16],en[8]);
bufif1 (Y[8],X[17],en[9]);
bufif1 (Y[8],X[18],en[10]);
bufif1 (Y[8],X[19],en[11]);
bufif1 (Y[8],X[20],en[12]);
bufif1 (Y[8],X[21],en[13]);
bufif1 (Y[8],X[22],en[14]);
bufif1 (Y[8],X[23],en[15]);

bufif1 (Y[9],X[9],en[0]);
bufif1 (Y[9],X[10],en[1]);
bufif1 (Y[9],X[11],en[2]);
bufif1 (Y[9],X[12],en[3]);
bufif1 (Y[9],X[13],en[4]);
bufif1 (Y[9],X[14],en[5]);
bufif1 (Y[9],X[15],en[6]);
bufif1 (Y[9],X[16],en[7]);
bufif1 (Y[9],X[17],en[8]);
bufif1 (Y[9],X[18],en[9]);
bufif1 (Y[9],X[19],en[10]);
bufif1 (Y[9],X[20],en[11]);
bufif1 (Y[9],X[21],en[12]);
bufif1 (Y[9],X[22],en[13]);
bufif1 (Y[9],X[23],en[14]);


bufif1 (Y[10],X[10],en[0]);
bufif1 (Y[10],X[11],en[1]);
bufif1 (Y[10],X[12],en[2]);
bufif1 (Y[10],X[13],en[3]);
bufif1 (Y[10],X[14],en[4]);
bufif1 (Y[10],X[15],en[5]);
bufif1 (Y[10],X[16],en[6]);
bufif1 (Y[10],X[17],en[7]);
bufif1 (Y[10],X[18],en[8]);
bufif1 (Y[10],X[19],en[9]);
bufif1 (Y[10],X[20],en[10]);
bufif1 (Y[10],X[21],en[11]);
bufif1 (Y[10],X[22],en[12]);
bufif1 (Y[10],X[23],en[13]);

bufif1 (Y[11],X[11],en[0]);
bufif1 (Y[11],X[12],en[1]);
bufif1 (Y[11],X[13],en[2]);
bufif1 (Y[11],X[14],en[3]);
bufif1 (Y[11],X[15],en[4]);
bufif1 (Y[11],X[16],en[5]);
bufif1 (Y[11],X[17],en[6]);
bufif1 (Y[11],X[18],en[7]);
bufif1 (Y[11],X[19],en[8]);
bufif1 (Y[11],X[20],en[9]);
bufif1 (Y[11],X[21],en[10]);
bufif1 (Y[11],X[22],en[11]);
bufif1 (Y[11],X[23],en[12]);

bufif1 (Y[12],X[12],en[0]);
bufif1 (Y[12],X[13],en[1]);
bufif1 (Y[12],X[14],en[2]);
bufif1 (Y[12],X[15],en[3]);
bufif1 (Y[12],X[16],en[4]);
bufif1 (Y[12],X[17],en[5]);
bufif1 (Y[12],X[18],en[6]);
bufif1 (Y[12],X[19],en[7]);
bufif1 (Y[12],X[20],en[8]);
bufif1 (Y[12],X[21],en[9]);
bufif1 (Y[12],X[22],en[10]);
bufif1 (Y[12],X[23],en[11]);

bufif1 (Y[13],X[13],en[0]);
bufif1 (Y[13],X[14],en[1]);
bufif1 (Y[13],X[15],en[2]);
bufif1 (Y[13],X[16],en[3]);
bufif1 (Y[13],X[17],en[4]);
bufif1 (Y[13],X[18],en[5]);
bufif1 (Y[13],X[19],en[6]);
bufif1 (Y[13],X[20],en[7]);
bufif1 (Y[13],X[21],en[8]);
bufif1 (Y[13],X[22],en[9]);
bufif1 (Y[13],X[23],en[10]);

bufif1 (Y[14],X[14],en[0]);
bufif1 (Y[14],X[15],en[1]);
bufif1 (Y[14],X[16],en[2]);
bufif1 (Y[14],X[17],en[3]);
bufif1 (Y[14],X[18],en[4]);
bufif1 (Y[14],X[19],en[5]);
bufif1 (Y[14],X[20],en[6]);
bufif1 (Y[14],X[21],en[7]);
bufif1 (Y[14],X[22],en[8]);
bufif1 (Y[14],X[23],en[9]);

bufif1 (Y[15],X[15],en[0]);
bufif1 (Y[15],X[16],en[1]);
bufif1 (Y[15],X[17],en[2]);
bufif1 (Y[15],X[18],en[3]);
bufif1 (Y[15],X[19],en[4]);
bufif1 (Y[15],X[20],en[5]);
bufif1 (Y[15],X[21],en[6]);
bufif1 (Y[15],X[22],en[7]);
bufif1 (Y[15],X[23],en[8]);

bufif1 (Y[16],X[16],en[0]);
bufif1 (Y[16],X[17],en[1]);
bufif1 (Y[16],X[18],en[2]);
bufif1 (Y[16],X[19],en[3]);
bufif1 (Y[16],X[20],en[4]);
bufif1 (Y[16],X[21],en[5]);
bufif1 (Y[16],X[22],en[6]);
bufif1 (Y[16],X[23],en[7]);

bufif1 (Y[17],X[17],en[0]);
bufif1 (Y[17],X[18],en[1]);
bufif1 (Y[17],X[19],en[2]);
bufif1 (Y[17],X[20],en[3]);
bufif1 (Y[17],X[21],en[4]);
bufif1 (Y[17],X[22],en[5]);
bufif1 (Y[17],X[23],en[6]);

bufif1 (Y[18],X[18],en[0]);
bufif1 (Y[18],X[19],en[1]);
bufif1 (Y[18],X[20],en[2]);
bufif1 (Y[18],X[21],en[3]);
bufif1 (Y[18],X[22],en[4]);
bufif1 (Y[18],X[23],en[5]);

bufif1 (Y[19],X[19],en[0]);
bufif1 (Y[19],X[20],en[1]);
bufif1 (Y[19],X[21],en[2]);
bufif1 (Y[19],X[22],en[3]);
bufif1 (Y[19],X[23],en[4]);

bufif1 (Y[20],X[20],en[0]);
bufif1 (Y[20],X[21],en[1]);
bufif1 (Y[20],X[22],en[2]);
bufif1 (Y[20],X[23],en[3]);

bufif1 (Y[21],X[21],en[0]);
bufif1 (Y[21],X[22],en[1]);
bufif1 (Y[21],X[23],en[2]);

bufif1 (Y[22],X[22],en[0]);
bufif1 (Y[22],X[23],en[1]);

bufif1 (Y[23],X[23],en[0]);

bufif1 (Y[0],0,en[24]);
or(en23,en[24],en[23]);
bufif1 (Y[1],0,en23);
or(en22,en23,en[22]);
bufif1 (Y[2],0,en22);
or(en21,en22,en[21]);
bufif1 (Y[3],0,en21);
or(en20,en21,en[20]);
bufif1 (Y[4],0,en20);
or(en19,en20,en[19]);
bufif1 (Y[5],0,en19);
or(en18,en19,en[18]);
bufif1 (Y[6],0,en18);
or(en17,en18,en[17]);
bufif1 (Y[7],0,en17);
or(en16,en17,en[16]);
bufif1 (Y[8],0,en16);
or(en15,en16,en[15]);
bufif1 (Y[9],0,en15);
or(en14,en15,en[14]);
bufif1 (Y[10],0,en14);
or(en13,en14,en[13]);
bufif1 (Y[11],0,en13);
or(en12,en13,en[12]);
bufif1 (Y[12],0,en12);
or(en11,en12,en[11]);
bufif1 (Y[13],0,en11);
or(en10,en11,en[10]);
bufif1 (Y[14],0,en10);
or(en9,en10,en[9]);
bufif1 (Y[15],0,en9);
or(en8,en9,en[8]);
bufif1 (Y[16],0,en8);
or(en7,en8,en[7]);
bufif1 (Y[17],0,en7);
or(en6,en7,en[6]);
bufif1 (Y[18],0,en6);
or(en5,en6,en[5]);
bufif1 (Y[19],0,en5);
or(en4,en5,en[4]);
bufif1 (Y[20],0,en4);
or(en3,en4,en[3]);
bufif1 (Y[21],0,en3);
or(en2,en3,en[2]);
bufif1 (Y[22],0,en2);
or(en1,en2,en[1]);
bufif1 (Y[23],0,en1);

endmodule 
