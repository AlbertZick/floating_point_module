module WallaceTree(a,b,c,d,e,f,g,h,i,j,k,l,m,out);
	input [25:0] a,b,c,d,e,f,g,h,i,j,k,l,m;
	output [47:0] out;

//Stage 0
HalfAdder H00(a[02],b[00],X2l,X2h);
HalfAdder H01(a[03],b[01],X3l,X3h);
FullAdder F0000(a[04],b[02],c[00],X4l,X4h);
FullAdder F0001(a[05],b[03],c[01],X5l,X5h);
FullAdder F0002(a[06],b[04],c[02],X6l,X6h);
FullAdder F0003(a[07],b[05],c[03],X7l,X7h);
FullAdder F0004(a[08],b[06],c[04],X8l,X8h);
FullAdder F0005(a[09],b[07],c[05],X9l,X9h);
FullAdder F0006(a[10],b[08],c[06],X10l,X10h);
FullAdder F0007(a[11],b[09],c[07],X11l,X11h);
FullAdder F0008(a[12],b[10],c[08],X12l,X12h);
FullAdder F0009(a[13],b[11],c[09],X13l,X13h);
FullAdder F0010(a[14],b[12],c[10],X14l,X14h);
FullAdder F0011(a[15],b[13],c[11],X15l,X15h);
FullAdder F0012(a[16],b[14],c[12],X16l,X16h);
FullAdder F0013(a[17],b[15],c[13],X17l,X17h);
FullAdder F0014(a[18],b[16],c[14],X18l,X18h);
FullAdder F0015(a[19],b[17],c[15],X19l,X19h);
FullAdder F0016(a[20],b[18],c[16],X20l,X20h);
FullAdder F0017(a[21],b[19],c[17],X21l,X21h);
FullAdder F0018(a[22],b[20],c[18],X22l,X22h);
FullAdder F0019(a[23],b[21],c[19],X23l,X23h);
FullAdder F0020(a[24],b[22],c[20],X24l,X24h);
FullAdder F0021(a[25],b[23],c[21],X25l,X25h);
FullAdder F0022(a[25],b[24],c[22],X26l,X26h);
FullAdder F0023(a[25],b[25],c[23],X27l,X27h);
FullAdder F0024(a[25],b[25],c[24],X28l,X28h);
FullAdder F0025(a[25],b[25],c[25],X29l,X29h);
FullAdder F0026(a[25],b[25],c[25],X30l,X30h);
FullAdder F0027(a[25],b[25],c[25],X31l,X31h);
FullAdder F0028(a[25],b[25],c[25],X32l,X32h);
FullAdder F0029(a[25],b[25],c[25],X33l,X33h);
FullAdder F0030(a[25],b[25],c[25],X34l,X34h);
FullAdder F0031(a[25],b[25],c[25],X35l,X35h);
FullAdder F0032(a[25],b[25],c[25],X36l,X36h);
FullAdder F0033(a[25],b[25],c[25],X37l,X37h);
FullAdder F0034(a[25],b[25],c[25],X38l,X38h);
FullAdder F0035(a[25],b[25],c[25],X39l,X39h);
FullAdder F0036(a[25],b[25],c[25],X40l,X40h);
FullAdder F0037(a[25],b[25],c[25],X41l,X41h);
FullAdder F0038(a[25],b[25],c[25],X42l,X42h);
FullAdder F0039(a[25],b[25],c[25],X43l,X43h);
FullAdder F0040(a[25],b[25],c[25],X44l,X44h);
FullAdder F0041(a[25],b[25],c[25],X45l,X45h);
FullAdder F0042(a[25],b[25],c[25],X46l,X46h);
FullAdder F0043(a[25],b[25],c[25],X47l,X47h);
FullAdder F0044(a[25],b[25],c[25],X48l,X48h);
FullAdder F0045(a[25],b[25],c[25],X49l,X49h);

HalfAdder H02(d[02],d[00],Y8l,Y8h);
HalfAdder H03(d[03],d[01],Y9l,Y9h);
FullAdder F0046(d[04],e[02],f[00],Y10l,Y10h);
FullAdder F0047(d[05],e[03],f[01],Y11l,Y11h);
FullAdder F0048(d[06],e[04],f[02],Y12l,Y12h);
FullAdder F0049(d[07],e[05],f[03],Y13l,Y13h);
FullAdder F0050(d[08],e[06],f[04],Y14l,Y14h);
FullAdder F0051(d[09],e[07],f[05],Y15l,Y15h);
FullAdder F0052(d[10],e[08],f[06],Y16l,Y16h);
FullAdder F0053(d[11],e[09],f[07],Y17l,Y17h);
FullAdder F0054(d[12],e[10],f[08],Y18l,Y18h);
FullAdder F0055(d[13],e[11],f[09],Y19l,Y19h);
FullAdder F0056(d[14],e[12],f[10],Y20l,Y20h);
FullAdder F0057(d[15],e[13],f[11],Y21l,Y21h);
FullAdder F0058(d[16],e[14],f[12],Y22l,Y22h);
FullAdder F0059(d[17],e[15],f[13],Y23l,Y23h);
FullAdder F0060(d[18],e[16],f[14],Y24l,Y24h);
FullAdder F0061(d[19],e[17],f[15],Y25l,Y25h);
FullAdder F0062(d[20],e[18],f[16],Y26l,Y26h);
FullAdder F0063(d[21],e[19],f[17],Y27l,Y27h);
FullAdder F0064(d[22],e[20],f[18],Y28l,Y28h);
FullAdder F0065(d[23],e[21],f[19],Y29l,Y29h);
FullAdder F0066(d[24],e[22],f[20],Y30l,Y30h);
FullAdder F0067(d[25],e[23],f[21],Y31l,Y31h);
FullAdder F0068(d[25],e[24],f[22],Y32l,Y32h);
FullAdder F0069(d[25],e[25],f[23],Y33l,Y33h);
FullAdder F0070(d[25],e[25],f[24],Y34l,Y34h);
FullAdder F0071(d[25],e[25],f[25],Y35l,Y35h);
FullAdder F0072(d[25],e[25],f[25],Y36l,Y36h);
FullAdder F0073(d[25],e[25],f[25],Y37l,Y37h);
FullAdder F0074(d[25],e[25],f[25],Y38l,Y38h);
FullAdder F0075(d[25],e[25],f[25],Y39l,Y39h);
FullAdder F0076(d[25],e[25],f[25],Y40l,Y40h);
FullAdder F0077(d[25],e[25],f[25],Y41l,Y41h);
FullAdder F0078(d[25],e[25],f[25],Y42l,Y42h);
FullAdder F0079(d[25],e[25],f[25],Y43l,Y43h);
FullAdder F0080(d[25],e[25],f[25],Y44l,Y44h);
FullAdder F0081(d[25],e[25],f[25],Y45l,Y45h);
FullAdder F0082(d[25],e[25],f[25],Y46l,Y46h);
FullAdder F0083(d[25],e[25],f[25],Y47l,Y47h);
FullAdder F0084(d[25],e[25],f[25],Y48l,Y48h);
FullAdder F0085(d[25],e[25],f[25],Y49l,Y49h);

HalfAdder H04(g[02],h[00],Z14l,Z14h);
HalfAdder H05(g[03],h[01],Z15l,Z15h);
FullAdder F0086(g[04],h[02],i[00],Z16l,Z16h);
FullAdder F0087(g[05],h[03],i[01],Z17l,Z17h);
FullAdder F0088(g[06],h[04],i[02],Z18l,Z18h);
FullAdder F0089(g[07],h[05],i[03],Z19l,Z19h);
FullAdder F0090(g[08],h[06],i[04],Z20l,Z20h);
FullAdder F0091(g[09],h[07],i[05],Z21l,Z21h);
FullAdder F0092(g[10],h[08],i[06],Z22l,Z22h);
FullAdder F0093(g[11],h[09],i[07],Z23l,Z23h);
FullAdder F0094(g[12],h[10],i[08],Z24l,Z24h);
FullAdder F0095(g[13],h[11],i[09],Z25l,Z25h);
FullAdder F0096(g[14],h[12],i[10],Z26l,Z26h);
FullAdder F0097(g[15],h[13],i[11],Z27l,Z27h);
FullAdder F0098(g[16],h[14],i[12],Z28l,Z28h);
FullAdder F0099(g[17],h[15],i[13],Z29l,Z29h);
FullAdder F0100(g[18],h[16],i[14],Z30l,Z30h);
FullAdder F0101(g[19],h[17],i[15],Z31l,Z31h);
FullAdder F0102(g[20],h[18],i[16],Z32l,Z32h);
FullAdder F0103(g[21],h[19],i[17],Z33l,Z33h);
FullAdder F0104(g[22],h[20],i[18],Z34l,Z34h);
FullAdder F0105(g[23],h[21],i[19],Z35l,Z35h);
FullAdder F0106(g[24],h[22],i[20],Z36l,Z36h);
FullAdder F0107(g[25],h[23],i[21],Z37l,Z37h);
FullAdder F0108(g[25],h[24],i[22],Z38l,Z38h);
FullAdder F0109(g[25],h[25],i[23],Z39l,Z39h);
FullAdder F0110(g[25],h[25],i[24],Z40l,Z40h);
FullAdder F0111(g[25],h[25],i[25],Z41l,Z41h);
FullAdder F0112(g[25],h[25],i[25],Z42l,Z42h);
FullAdder F0113(g[25],h[25],i[25],Z43l,Z43h);
FullAdder F0114(g[25],h[25],i[25],Z44l,Z44h);
FullAdder F0115(g[25],h[25],i[25],Z45l,Z45h);
FullAdder F0116(g[25],h[25],i[25],Z46l,Z46h);
FullAdder F0117(g[25],h[25],i[25],Z47l,Z47h);
FullAdder F0118(g[25],h[25],i[25],Z48l,Z48h);
FullAdder F0119(g[25],h[25],i[25],Z49l,Z49h);

HalfAdder H06(j[02],k[00],T20l,T20h);
HalfAdder H07(j[03],k[01],T21l,T21h);
FullAdder F0120(j[04],k[02],l[00],T22l,T22h);
FullAdder F0121(j[05],k[03],l[01],T23l,T23h);
FullAdder F0122(j[06],k[04],l[02],T24l,T24h);
FullAdder F0123(j[07],k[05],l[03],T25l,T25h);
FullAdder F0124(j[08],k[06],l[04],T26l,T26h);
FullAdder F0125(j[09],k[07],l[05],T27l,T27h);
FullAdder F0126(j[10],k[08],l[06],T28l,T28h);
FullAdder F0127(j[11],k[09],l[07],T29l,T29h);
FullAdder F0128(j[12],k[10],l[08],T30l,T30h);
FullAdder F0129(j[13],k[11],l[09],T31l,T31h);
FullAdder F0130(j[14],k[12],l[10],T32l,T32h);
FullAdder F0131(j[15],k[13],l[11],T33l,T33h);
FullAdder F0132(j[16],k[14],l[12],T34l,T34h);
FullAdder F0133(j[17],k[15],l[13],T35l,T35h);
FullAdder F0134(j[18],k[16],l[14],T36l,T36h);
FullAdder F0135(j[19],k[17],l[15],T37l,T37h);
FullAdder F0136(j[20],k[18],l[16],T38l,T38h);
FullAdder F0137(j[21],k[19],l[17],T39l,T39h);
FullAdder F0138(j[22],k[20],l[18],T40l,T40h);
FullAdder F0139(j[23],k[21],l[19],T41l,T41h);
FullAdder F0140(j[24],k[22],l[20],T42l,T42h);
FullAdder F0141(j[25],k[23],l[21],T43l,T43h);
FullAdder F0142(j[25],k[24],l[22],T44l,T44h);
FullAdder F0143(j[25],k[25],l[23],T45l,T45h);
FullAdder F0144(j[25],k[25],l[24],T46l,T46h);
FullAdder F0145(j[25],k[25],l[25],T47l,T47h);
FullAdder F0146(j[25],k[25],l[25],T48l,T48h);
FullAdder F0147(j[25],k[25],l[25],T49l,T49h);



//Stage 1
HalfAdder H10(X2h,X3l,XX3l,XX3h);
HalfAdder H11(X3h,X4l,XX4l,XX4h);
HalfAdder H12(X4h,X5l,XX5l,XX5h);
FullAdder F101(X5h,X6l,d[0],XX6l,XX6h);
FullAdder F102(X6h,X7l,d[1],XX7l,XX7h);
FullAdder F103(X7h,X8l,Y8l,XX8l,XX8h);
FullAdder F104(X8h,Y8h,X9l,XX9l,XX9h);
FullAdder F105(X9h,Y9h,X10l,XX10l,XX10h);
FullAdder F106(X10h,Y10h,X11l,XX11l,XX11h);
FullAdder F107(X11h,Y11h,X12l,XX12l,XX12h);
FullAdder F108(X12h,Y12h,X13l,XX13l,XX13h);
FullAdder F109(X13h,Y13h,X14l,XX14l,XX14h);
FullAdder F110(X14h,Y14h,Z14h,XX15l,XX15h);
FullAdder F111(X15h,Y15h,Z15h,XX16l,XX16h);
FullAdder F112(X16h,Y16h,Z16h,XX17l,XX17h);
FullAdder F113(X17h,Y17h,Z17h,XX18l,XX18h);
FullAdder F114(X18h,Y18h,Z18h,XX19l,XX19h);
FullAdder F115(X19h,Y19h,Z19h,XX20l,XX20h);
FullAdder F116(X20h,Y20h,Z20h,XX21l,XX21h);
FullAdder F117(X21h,Y21h,Z21h,XX22l,XX22h);
FullAdder F118(X22h,Y22h,Z22h,XX23l,XX23h);
FullAdder F119(X23h,Y23h,Z23h,XX24l,XX24h);
FullAdder F120(X24h,Y24h,Z24h,XX25l,XX25h);
FullAdder F121(X25h,Y25h,Z25h,XX26l,XX26h);
FullAdder F122(X26h,Y26h,Z26h,XX27l,XX27h);
FullAdder F123(X27h,Y27h,Z27h,XX28l,XX28h);
FullAdder F124(X28h,Y28h,Z28h,XX29l,XX29h);
FullAdder F125(X29h,Y29h,Z29h,XX30l,XX30h);
FullAdder F126(X30h,Y30h,Z30h,XX31l,XX31h);
FullAdder F127(X31h,Y31h,Z31h,XX32l,XX32h);
FullAdder F128(X32h,Y32h,Z32h,XX33l,XX33h);
FullAdder F129(X33h,Y33h,Z33h,XX34l,XX34h);
FullAdder F130(X34h,Y34h,Z34h,XX35l,XX35h);
FullAdder F131(X35h,Y35h,Z35h,XX36l,XX36h);
FullAdder F132(X36h,Y36h,Z36h,XX37l,XX37h);
FullAdder F133(X37h,Y37h,Z37h,XX38l,XX38h);
FullAdder F134(X38h,Y38h,Z38h,XX39l,XX39h);
FullAdder F135(X39h,Y39h,Z39h,XX40l,XX40h);
FullAdder F136(X40h,Y40h,Z40h,XX41l,XX41h);
FullAdder F137(X41h,Y41h,Z41h,XX42l,XX42h);
FullAdder F138(X42h,Y42h,Z42h,XX43l,XX43h);
FullAdder F139(X43h,Y43h,Z43h,XX44l,XX44h);
FullAdder F140(X44h,Y44h,Z44h,XX45l,XX45h);
FullAdder F141(X45h,Y45h,Z45h,XX46l,XX46h);
FullAdder F142(X46h,Y46h,Z46h,XX47l,XX47h);
FullAdder F143(X47h,Y47h,Z47h,XX48l,XX48h);
FullAdder F144(X48h,Y48h,Z48h,XX49l,XX49h);

HalfAdder H13(Y12l,g[0],YY12l,YY12h);
HalfAdder H14(Y13l,g[1],YY13l,YY13h);
HalfAdder H15(Y14l,Z14l,YY14l,YY14h);
FullAdder F146(X15l,Y15l,Z15l,YY15l,YY15h);
FullAdder F147(X16l,Y16l,Z16l,YY16l,YY16h);
FullAdder F148(X17l,Y17l,Z17l,YY17l,YY17h);
FullAdder F149(X18l,Y18l,Z18l,YY18l,YY18h);
FullAdder F150(X19l,Y19l,Z19l,YY19l,YY19h);
FullAdder F151(X20l,Y20l,Z20l,YY20l,YY20h);
FullAdder F152(T20h,X21l,Y21l,YY21l,YY21h);
FullAdder F153(T21h,X22l,Y22l,YY22l,YY22h);
FullAdder F154(T22h,X23l,Y23l,YY23l,YY23h);
FullAdder F155(T23h,X24l,Y24l,YY24l,YY24h);
FullAdder F156(T24h,X25l,Y25l,YY25l,YY25h);
FullAdder F157(T25h,X26l,Y26l,YY26l,YY26h);
FullAdder F158(T26h,X27l,Y27l,YY27l,YY27h);
FullAdder F159(T27h,X28l,Y28l,YY28l,YY28h);
FullAdder F160(T28h,X29l,Y29l,YY29l,YY29h);
FullAdder F161(T29h,X30l,Y30l,YY30l,YY30h);
FullAdder F162(T30h,X31l,Y31l,YY31l,YY31h);
FullAdder F163(T31h,X32l,Y32l,YY32l,YY32h);
FullAdder F164(T32h,X33l,Y33l,YY33l,YY33h);
FullAdder F165(T33h,X34l,Y34l,YY34l,YY34h);
FullAdder F166(T34h,X35l,Y35l,YY35l,YY35h);
FullAdder F167(T35h,X36l,Y36l,YY36l,YY36h);
FullAdder F168(T36h,X37l,Y37l,YY37l,YY37h);
FullAdder F169(T37h,X38l,Y38l,YY38l,YY38h);
FullAdder F170(T38h,X39l,Y39l,YY39l,YY39h);
FullAdder F171(T39h,X40l,Y40l,YY40l,YY40h);
FullAdder F172(T40h,X41l,Y41l,YY41l,YY41h);
FullAdder F173(T41h,X42l,Y42l,YY42l,YY42h);
FullAdder F174(T42h,X43l,Y43l,YY43l,YY43h);
FullAdder F175(T43h,X44l,Y44l,YY44l,YY44h);
FullAdder F176(T44h,X45l,Y45l,YY45l,YY45h);
FullAdder F177(T45h,X46l,Y46l,YY46l,YY46h);
FullAdder F178(T46h,X47l,Y47l,YY47l,YY47h);
FullAdder F179(T47h,X48l,Y48l,YY48l,YY48h);
FullAdder F180(T48h,X49l,Y49l,YY49l,YY49h);

HalfAdder H16(Z21l,T21l,ZZ21l,ZZ21h);
HalfAdder H17(Z22l,T22l,ZZ22l,ZZ22h);
HalfAdder H18(Z23l,T23l,ZZ23l,ZZ23h);
FullAdder F181(Z24l,T24l,m[00],ZZ24l,ZZ24h);
FullAdder F182(Z25l,T25l,m[01],ZZ25l,ZZ25h);
FullAdder F183(Z26l,T26l,m[02],ZZ26l,ZZ26h);
FullAdder F184(Z27l,T27l,m[03],ZZ27l,ZZ27h);
FullAdder F185(Z28l,T28l,m[04],ZZ28l,ZZ28h);
FullAdder F186(Z29l,T29l,m[05],ZZ29l,ZZ29h);
FullAdder F187(Z30l,T30l,m[06],ZZ30l,ZZ30h);
FullAdder F188(Z31l,T31l,m[07],ZZ31l,ZZ31h);
FullAdder F189(Z32l,T32l,m[08],ZZ32l,ZZ32h);
FullAdder F190(Z33l,T33l,m[09],ZZ33l,ZZ33h);
FullAdder F191(Z34l,T34l,m[10],ZZ34l,ZZ34h);
FullAdder F192(Z35l,T35l,m[11],ZZ35l,ZZ35h);
FullAdder F193(Z36l,T36l,m[12],ZZ36l,ZZ36h);
FullAdder F194(Z37l,T37l,m[13],ZZ37l,ZZ37h);
FullAdder F195(Z38l,T38l,m[14],ZZ38l,ZZ38h);
FullAdder F196(Z39l,T39l,m[15],ZZ39l,ZZ39h);
FullAdder F197(Z40l,T40l,m[16],ZZ40l,ZZ40h);
FullAdder F198(Z41l,T41l,m[17],ZZ41l,ZZ41h);
FullAdder F199(Z42l,T42l,m[18],ZZ42l,ZZ42h);
FullAdder F1101(Z43l,T43l,m[19],ZZ43l,ZZ43h);
FullAdder F1102(Z44l,T44l,m[20],ZZ44l,ZZ44h);
FullAdder F1103(Z45l,T45l,m[21],ZZ45l,ZZ45h);
FullAdder F1104(Z46l,T46l,m[22],ZZ46l,ZZ46h);
FullAdder F1105(Z47l,T47l,m[23],ZZ47l,ZZ47h);
FullAdder F1106(Z48l,T48l,m[24],ZZ48l,ZZ48h);
FullAdder F1107(Z49l,T49l,m[25],ZZ49l,ZZ49h);




//Stage 2
HalfAdder H20(XX3h,XX4l,XXX4l,XXX4h);
HalfAdder H21(XX4h,XX5l,XXX5l,XXX5h);
HalfAdder H22(XX5h,XX6l,XXX6l,XXX6h);
HalfAdder H23(XX6h,XX7l,XXX7l,XXX7h);
HalfAdder H24(XX7h,XX8l,XXX8l,XXX8h);
FullAdder F200(XX8h,XX9l,Y9l,XXX9l,XXX9h);
FullAdder F201(XX9h,XX10l,Y10l,XXX10l,XXX10h);
FullAdder F202(XX10h,XX11l,Y11l,XXX11l,XXX11h);
FullAdder F203(XX11h,XX12l,YY12l,XXX12l,XXX12h);
FullAdder F204(XX12h,YY12h,XX13l,XXX13l,XXX13h);
FullAdder F205(XX13h,YY13h,XX14l,XXX14l,XXX14h);
FullAdder F206(XX14h,YY14h,XX15l,XXX15l,XXX15h);
FullAdder F207(XX15h,YY15h,XX16l,XXX16l,XXX16h);
FullAdder F208(XX16h,YY16h,XX17l,XXX17l,XXX17h);
FullAdder F209(XX17h,YY17h,XX18l,XXX18l,XXX18h);
FullAdder F210(XX18h,YY18h,XX19l,XXX19l,XXX19h);
FullAdder F211(XX19h,YY19h,XX20l,XXX20l,XXX20h);
FullAdder F212(XX20h,YY20h,XX21l,XXX21l,XXX21h);
FullAdder F213(XX21h,YY21h,ZZ21h,XXX22l,XXX22h);
FullAdder F214(XX22h,YY22h,ZZ22h,XXX23l,XXX23h);
FullAdder F215(XX23h,YY23h,ZZ23h,XXX24l,XXX24h);
FullAdder F216(XX24h,YY24h,ZZ24h,XXX25l,XXX25h);
FullAdder F217(XX25h,YY25h,ZZ25h,XXX26l,XXX26h);
FullAdder F218(XX26h,YY26h,ZZ26h,XXX27l,XXX27h);
FullAdder F219(XX27h,YY27h,ZZ27h,XXX28l,XXX28h);
FullAdder F220(XX28h,YY28h,ZZ28h,XXX29l,XXX29h);
FullAdder F221(XX29h,YY29h,ZZ29h,XXX30l,XXX30h);
FullAdder F222(XX30h,YY30h,ZZ30h,XXX31l,XXX31h);
FullAdder F223(XX31h,YY31h,ZZ31h,XXX32l,XXX32h);
FullAdder F224(XX32h,YY32h,ZZ32h,XXX33l,XXX33h);
FullAdder F225(XX33h,YY33h,ZZ33h,XXX34l,XXX34h);
FullAdder F226(XX34h,YY34h,ZZ34h,XXX35l,XXX35h);
FullAdder F227(XX35h,YY35h,ZZ35h,XXX36l,XXX36h);
FullAdder F228(XX36h,YY36h,ZZ36h,XXX37l,XXX37h);
FullAdder F229(XX37h,YY37h,ZZ37h,XXX38l,XXX38h);
FullAdder F230(XX38h,YY38h,ZZ38h,XXX39l,XXX39h);
FullAdder F231(XX39h,YY39h,ZZ39h,XXX40l,XXX40h);
FullAdder F232(XX40h,YY40h,ZZ40h,XXX41l,XXX41h);
FullAdder F233(XX41h,YY41h,ZZ41h,XXX42l,XXX42h);
FullAdder F234(XX42h,YY42h,ZZ42h,XXX43l,XXX43h);
FullAdder F235(XX43h,YY43h,ZZ43h,XXX44l,XXX44h);
FullAdder F236(XX44h,YY44h,ZZ44h,XXX45l,XXX45h);
FullAdder F237(XX45h,YY45h,ZZ45h,XXX46l,XXX46h);
FullAdder F238(XX46h,YY46h,ZZ46h,XXX47l,XXX47h);
FullAdder F239(XX47h,YY47h,ZZ47h,XXX48l,XXX48h);
FullAdder F240(XX48h,YY48h,ZZ48h,XXX49l,XXX49h);

HalfAdder H25(YY18l,j[0],YYY18l,YYY18h);
HalfAdder H26(YY19l,j[1],YYY19l,YYY19h);
HalfAdder H27(YY20l,T20l,YYY20l,YYY20h);
HalfAdder H28(YY21l,ZZ21l,YYY21l,YYY21h);
FullAdder F241(XX22l,YY22l,ZZ22l,YYY22l,YYY22h);
FullAdder F242(XX23l,YY23l,ZZ23l,YYY23l,YYY23h);
FullAdder F243(XX24l,YY24l,ZZ24l,YYY24l,YYY24h);
FullAdder F244(XX25l,YY25l,ZZ25l,YYY25l,YYY25h);
FullAdder F245(XX26l,YY26l,ZZ26l,YYY26l,YYY26h);
FullAdder F246(XX27l,YY27l,ZZ27l,YYY27l,YYY27h);
FullAdder F247(XX28l,YY28l,ZZ28l,YYY28l,YYY28h);
FullAdder F248(XX29l,YY29l,ZZ29l,YYY29l,YYY29h);
FullAdder F249(XX30l,YY30l,ZZ30l,YYY30l,YYY30h);
FullAdder F250(XX31l,YY31l,ZZ31l,YYY31l,YYY31h);
FullAdder F251(XX32l,YY32l,ZZ32l,YYY32l,YYY32h);
FullAdder F252(XX33l,YY33l,ZZ33l,YYY33l,YYY33h);
FullAdder F253(XX34l,YY34l,ZZ34l,YYY34l,YYY34h);
FullAdder F254(XX35l,YY35l,ZZ35l,YYY35l,YYY35h);
FullAdder F255(XX36l,YY36l,ZZ36l,YYY36l,YYY36h);
FullAdder F256(XX37l,YY37l,ZZ37l,YYY37l,YYY37h);
FullAdder F257(XX38l,YY38l,ZZ38l,YYY38l,YYY38h);
FullAdder F258(XX39l,YY39l,ZZ39l,YYY39l,YYY39h);
FullAdder F259(XX40l,YY40l,ZZ40l,YYY40l,YYY40h);
FullAdder F260(XX41l,YY41l,ZZ41l,YYY41l,YYY41h);
FullAdder F261(XX42l,YY42l,ZZ42l,YYY42l,YYY42h);
FullAdder F262(XX43l,YY43l,ZZ43l,YYY43l,YYY43h);
FullAdder F263(XX44l,YY44l,ZZ44l,YYY44l,YYY44h);
FullAdder F264(XX45l,YY45l,ZZ45l,YYY45l,YYY45h);
FullAdder F265(XX46l,YY46l,ZZ46l,YYY46l,YYY46h);
FullAdder F266(XX47l,YY47l,ZZ47l,YYY47l,YYY47h);
FullAdder F267(XX48l,YY48l,ZZ48l,YYY48l,YYY48h);
FullAdder F268(XX49l,YY49l,ZZ49l,YYY49l,YYY49h);



//Stage 3
HalfAdder H30(XXX4h,XXX5l,M5l,M5h);
HalfAdder H31(XXX5h,XXX6l,M6l,M6h);
HalfAdder H32(XXX6h,XXX7l,M7l,M7h);
HalfAdder H33(XXX7h,XXX8l,M8l,M8h);
HalfAdder H34(XXX8h,XXX9l,M9l,M9h);
HalfAdder H35(XXX9h,XXX10l,M10l,M10h);
HalfAdder H36(XXX10h,XXX11l,M11l,M11h);
HalfAdder H37(XXX11h,XXX12l,M12l,M12h);
FullAdder F300(XXX12h,XXX13l,YY13l,M13l,M13h);
FullAdder F301(XXX13h,XXX14l,YY14l,M14l,M14h);
FullAdder F302(XXX14h,XXX15l,YY15l,M15l,M15h);
FullAdder F303(XXX15h,XXX16l,YY16l,M16l,M16h);
FullAdder F304(XXX16h,XXX17l,YY17l,M17l,M17h);
FullAdder F305(XXX17h,XXX18l,YYY18l,M18l,M18h);
FullAdder F306(XXX18h,YYY18h,XXX19l,M19l,M19h);
FullAdder F307(XXX19h,YYY19h,XXX20l,M20l,M20h);
FullAdder F308(XXX20h,YYY20h,XXX21l,M21l,M21h);
FullAdder F309(XXX21h,YYY21h,XXX22l,M22l,M22h);
FullAdder F310(XXX22h,YYY22h,XXX23l,M23l,M23h);
FullAdder F311(XXX23h,YYY23h,XXX24l,M24l,M24h);
FullAdder F312(XXX24h,YYY24h,XXX25l,M25l,M25h);
FullAdder F313(XXX25h,YYY25h,XXX26l,M26l,M26h);
FullAdder F314(XXX26h,YYY26h,XXX27l,M27l,M27h);
FullAdder F315(XXX27h,YYY27h,XXX28l,M28l,M28h);
FullAdder F316(XXX28h,YYY28h,XXX29l,M29l,M29h);
FullAdder F317(XXX29h,YYY29h,XXX30l,M30l,M30h);
FullAdder F318(XXX30h,YYY30h,XXX31l,M31l,M31h);
FullAdder F319(XXX31h,YYY31h,XXX32l,M32l,M32h);
FullAdder F320(XXX32h,YYY32h,XXX33l,M33l,M33h);
FullAdder F321(XXX33h,YYY33h,XXX34l,M34l,M34h);
FullAdder F322(XXX34h,YYY34h,XXX35l,M35l,M35h);
FullAdder F323(XXX35h,YYY35h,XXX36l,M36l,M36h);
FullAdder F324(XXX36h,YYY36h,XXX37l,M37l,M37h);
FullAdder F325(XXX37h,YYY37h,XXX38l,M38l,M38h);
FullAdder F326(XXX38h,YYY38h,XXX39l,M39l,M39h);
FullAdder F327(XXX39h,YYY39h,XXX40l,M40l,M40h);
FullAdder F328(XXX40h,YYY40h,XXX41l,M41l,M41h);
FullAdder F329(XXX41h,YYY41h,XXX42l,M42l,M42h);
FullAdder F330(XXX42h,YYY42h,XXX43l,M43l,M43h);
FullAdder F331(XXX43h,YYY43h,XXX44l,M44l,M44h);
FullAdder F332(XXX44h,YYY44h,XXX45l,M45l,M45h);
FullAdder F333(XXX45h,YYY45h,XXX46l,M46l,M46h);
FullAdder F334(XXX46h,YYY46h,XXX47l,M47l,M47h);
FullAdder F335(XXX47h,YYY47h,XXX48l,M48l,M48h);
FullAdder F336(XXX48h,YYY48h,XXX49l,M49l,M49h);




//Stage 4
HalfAdder H400(M5h,M6l,MM6l,MM6h);
HalfAdder H401(M6h,M7l,MM7l,MM7h);
HalfAdder H402(M7h,M8l,MM8l,MM8h);
HalfAdder H403(M8h,M9l,MM9l,MM9h);
HalfAdder H404(M9h,M10l,MM10l,MM10h);
HalfAdder H405(M10h,M11l,MM11l,MM11h);
HalfAdder H406(M11h,M12l,MM12l,MM12h);
HalfAdder H407(M12h,M13l,MM13l,MM13h);
HalfAdder H408(M13h,M14l,MM14l,MM14h);
HalfAdder H409(M14h,M15l,MM15l,MM15h);
HalfAdder H410(M15h,M16l,MM16l,MM16h);
HalfAdder H411(M16h,M17l,MM17l,MM17h);
HalfAdder H412(M17h,M18l,MM18l,MM18h);
FullAdder F401(M18h,M19l,YYY19l,MM19l,MM19h);
FullAdder F402(M19h,M20l,YYY20l,MM20l,MM20h);
FullAdder F403(M20h,M21l,YYY21l,MM21l,MM21h);
FullAdder F404(M21h,M22l,YYY22l,MM22l,MM22h);
FullAdder F405(M22h,M23l,YYY23l,MM23l,MM23h);
FullAdder F406(M23h,M24l,YYY24l,MM24l,MM24h);
FullAdder F407(M24h,M25l,YYY25l,MM25l,MM25h);
FullAdder F408(M25h,M26l,YYY26l,MM26l,MM26h);
FullAdder F409(M26h,M27l,YYY27l,MM27l,MM27h);
FullAdder F410(M27h,M28l,YYY28l,MM28l,MM28h);
FullAdder F411(M28h,M29l,YYY29l,MM29l,MM29h);
FullAdder F412(M29h,M30l,YYY30l,MM30l,MM30h);
FullAdder F413(M30h,M31l,YYY31l,MM31l,MM31h);
FullAdder F414(M31h,M32l,YYY32l,MM32l,MM32h);
FullAdder F415(M32h,M33l,YYY33l,MM33l,MM33h);
FullAdder F416(M33h,M34l,YYY34l,MM34l,MM34h);
FullAdder F417(M34h,M35l,YYY35l,MM35l,MM35h);
FullAdder F418(M35h,M36l,YYY36l,MM36l,MM36h);
FullAdder F419(M36h,M37l,YYY37l,MM37l,MM37h);
FullAdder F420(M37h,M38l,YYY38l,MM38l,MM38h);
FullAdder F421(M38h,M39l,YYY39l,MM39l,MM39h);
FullAdder F422(M39h,M40l,YYY40l,MM40l,MM40h);
FullAdder F423(M40h,M41l,YYY41l,MM41l,MM41h);
FullAdder F424(M41h,M42l,YYY42l,MM42l,MM42h);
FullAdder F425(M42h,M43l,YYY43l,MM43l,MM43h);
FullAdder F426(M43h,M44l,YYY44l,MM44l,MM44h);
FullAdder F427(M44h,M45l,YYY45l,MM45l,MM45h);
FullAdder F428(M45h,M46l,YYY46l,MM46l,MM46h);
FullAdder F429(M46h,M47l,YYY47l,MM47l,MM47h);
FullAdder F430(M47h,M48l,YYY48l,MM48l,MM48h);
FullAdder F431(M48h,M49l,YYY49l,MM49l,MM49h);


//Final Stage
assign out[0]=a[0];
assign out[1]=a[1];
assign out[2]=X2l;
assign out[3]=XX3l;
assign out[4]=XXX4l;
assign out[5]=M5l;
assign out[6]=MM6l;
HalfAdder HF0(MM6h,MM7l,out[7],CR7);
FullAdder FF00(MM7h,MM8l,CR7,out[8],CR8);
FullAdder FF01(MM8h,MM9l,CR8,out[9],CR9);
FullAdder FF02(MM9h,MM10l,CR9,out[10],CR10);
FullAdder FF03(MM10h,MM11l,CR10,out[11],CR11);
FullAdder FF04(MM11h,MM12l,CR11,out[12],CR12);
FullAdder FF05(MM12h,MM13l,CR12,out[13],CR13);
FullAdder FF06(MM13h,MM14l,CR13,out[14],CR14);
FullAdder FF07(MM14h,MM15l,CR14,out[15],CR15);
FullAdder FF08(MM15h,MM16l,CR15,out[16],CR16);
FullAdder FF09(MM16h,MM17l,CR16,out[17],CR17);
FullAdder FF10(MM17h,MM18l,CR17,out[18],CR18);
FullAdder FF11(MM18h,MM19l,CR18,out[19],CR19);
FullAdder FF12(MM19h,MM20l,CR19,out[20],CR20);
FullAdder FF13(MM20h,MM21l,CR20,out[21],CR21);
FullAdder FF14(MM21h,MM22l,CR21,out[22],CR22);
FullAdder FF15(MM22h,MM23l,CR22,out[23],CR23);
FullAdder FF16(MM23h,MM24l,CR23,out[24],CR24);
FullAdder FF17(MM24h,MM25l,CR24,out[25],CR25);
FullAdder FF18(MM25h,MM26l,CR25,out[26],CR26);
FullAdder FF19(MM26h,MM27l,CR26,out[27],CR27);
FullAdder FF20(MM27h,MM28l,CR27,out[28],CR28);
FullAdder FF21(MM28h,MM29l,CR28,out[29],CR29);
FullAdder FF22(MM29h,MM30l,CR29,out[30],CR30);
FullAdder FF23(MM30h,MM31l,CR30,out[31],CR31);
FullAdder FF24(MM31h,MM32l,CR31,out[32],CR32);
FullAdder FF25(MM32h,MM33l,CR32,out[33],CR33);
FullAdder FF26(MM33h,MM34l,CR33,out[34],CR34);
FullAdder FF27(MM34h,MM35l,CR34,out[35],CR35);
FullAdder FF28(MM35h,MM36l,CR35,out[36],CR36);
FullAdder FF29(MM36h,MM37l,CR36,out[37],CR37);
FullAdder FF30(MM37h,MM38l,CR37,out[38],CR38);
FullAdder FF31(MM38h,MM39l,CR38,out[39],CR39);
FullAdder FF32(MM39h,MM40l,CR39,out[40],CR40);
FullAdder FF33(MM40h,MM41l,CR40,out[41],CR41);
FullAdder FF34(MM41h,MM42l,CR41,out[42],CR42);
FullAdder FF35(MM42h,MM43l,CR42,out[43],CR43);
FullAdder FF36(MM43h,MM44l,CR43,out[44],CR44);
FullAdder FF37(MM44h,MM45l,CR44,out[45],CR45);
FullAdder FF38(MM45h,MM46l,CR45,out[46],CR46);
FullAdder FF39(MM46h,MM47l,CR46,out[47],CR47);
// FullAdder FF40(MM47h,MM48l,CR47,out[48],CR48);
// FullAdder FF41(MM48h,MM49l,CR48,out[49],CR49);

endmodule