module Final_tb;
	reg clk,en,rst_n;
	reg [1:0] op; //00 = add; 01 = subtract; 10 = multiply; 11 = divide;
	reg [31:0] inA,inB;
	wire [31:0] out;
	wire finish;

	FloatingPointCalculator FPC(inA,inB,op,en,rst_n,clk,out,finish);

	initial begin
	clk = 0 ;
	en = 1 ;
	rst_n = 0 ;

	///////////////////////////////////////////////////////
	////              Add and subtract                 ////
	///////////////////////////////////////////////////////

	//Normal cases
	inA=32'b01000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//7.5 + 1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//7.5 + (-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b11000001000101110101110000101001; op=0;	//7.5 + (-9.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//(-7.5)+1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b01000001000101110101110000101001; op=0;	//(-7.5)+9.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//(-7.5)+(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//7.5 - 1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b01000001000101110101110000101001; op=1;	//7.5 - 9.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//7.5 - (-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//(-7.5)-1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//-7.5 - (-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b11000001000101110101110000101001; op=1;	//-7.5 - (-9.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b01000000111100000000000000000000; op=1;	//7.5 - 7.5
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b11000000111100000000000000000000; op=0;	//7.5 + (-7.5)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b01000000111100000000000000000000; op=0;	//-7.5 + 7.5
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b11000000111100000000000000000000; op=1;	//-7.5 - (-7.5)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	//Zero cases
	inA=32'b01000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=0; 	//7.5+0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=1; 	//7.5-0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=0; 	//-7.5+0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=1; 	//-7.5-0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//0+1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//0-1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//0+(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//0-(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;	//0+0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;	//0-0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	//Infinity cases
	inA=32'b01000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//7.5+inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//7.5-inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//7.5+(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//7.5-(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//-7.5+inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//-7.5-inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//-7.5+(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//-7.5-(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//inf+1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//inf-1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//inf+(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//inf-(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//-inf+1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//-inf-1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//-inf+(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//-inf-(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//inf+inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//inf-inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//inf+(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//inf-(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//-inf+inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//-inf-inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//-inf+(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//-inf-(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	//NaN cases
	inA=32'b01000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//7.5+NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//7.5+NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//-7.5+NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//-7.5-NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b00111111101110101110000101001000; op=0;	//NaN+1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b00111111101110101110000101001000; op=1;	//NaN-1.46
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b10111111101110101110000101001000; op=0;	//NaN+(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b10111111101110101110000101001000; op=1;	//NaN-(-1.46)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b01111111101010101010101010101010; op=0;	//NaN+NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b01111111101010101010101010101010; op=1;	//NaN-NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	//Crossover cases
	inA=32'b00000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//0+inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//0+inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//0+(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//0-(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;	//inf+0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;	//inf-0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;	//-inf+0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;	//-inf-0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//0+NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//0-NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b00000000000000000000000000000000; op=0;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b10000000000000000000000000000000; op=0;	//NaN+0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b00000000000000000000000000000000; op=1;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b10000000000000000000000000000000; op=1;	//NaN-0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//inf+NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//inf-NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//-inf+NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//-inf-NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b01111111100000000000000000000000; op=0;	//NaN+inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b01111111100000000000000000000000; op=1;	//NaN-inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b11111111100000000000000000000000; op=0;	//NaN+(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010;inB=32'b11111111100000000000000000000000; op=1;	//NaN-(-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;


	///////////////////////////////////////////////////////
	////                  Multiply                     ////
	///////////////////////////////////////////////////////
	op = 2'b10;
	//Normal cases
	inA=32'b00111111110000000000000000000000; inB=32'b01000010101110010101110000101001; //1.5 * 92.68
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111110000000000000000000000; inB=32'b11000010101110010101110000101001; //1.5 * (-92.68)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111110000000000000000000000; inB=32'b01000010101110010101110000101001; //-1.5 * 92.68
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111110000000000000000000000; inB=32'b11000010101110010101110000101001; //-1.5 * (-92.68)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	//Zero cases
	inA=32'b00000000000000000000000000000000; inB=32'b01000010101110010101110000101001; 
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01000010101110010101110000101001; //0 * 92.68
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b11000010101110010101110000101001; 
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b11000010101110010101110000101001; //0 * (-92.68)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111110000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111110000000000000000000000; inB=32'b10000000000000000000000000000000; //1.5 * 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111110000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111110000000000000000000000; inB=32'b10000000000000000000000000000000; //-1.5 * 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b10000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b10000000000000000000000000000000; //0 * 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	//Infinity cases
	inA=32'b01111111100000000000000000000000; inB=32'b01000010101110010101110000101001; //inf * 92.68
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01000010101110010101110000101001; //-inf * 92.68
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b11000010101110010101110000101001; //inf * (-92.68)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b11000010101110010101110000101001; //-inf * (-92.68)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111110000000000000000000000; inB=32'b01111111100000000000000000000000; //1.5 * inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111110000000000000000000000; inB=32'b11111111100000000000000000000000; //1.5 * (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111110000000000000000000000; inB=32'b01111111100000000000000000000000; //-1.5 * inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111110000000000000000000000; inB=32'b11111111100000000000000000000000; //-1.5 * (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	//inf * inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b11111111100000000000000000000000;	//inf * (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	//-inf * inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b11111111100000000000000000000000;	//-inf * (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	//NaN cases
	inA=32'b00111111110000000000000000000000; inB=32'b01111111101010101010101010101010; //1.5 * NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111110000000000000000000000; inB=32'b01111111101010101010101010101010; //-1.5 * NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b01000010101110010101110000101001; //NaN * 92.68
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b11000010101110010101110000101001; //NaN * (-92.68)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b01111111101010101010101010101010; //NaN * NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;	
	//Crossover cases
	inA=32'b00000000000000000000000000000000; inB=32'b01111111100000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01111111100000000000000000000000; //0 * inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b11111111100000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b11111111100000000000000000000000; //0 * (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b01111111101010101010101010101010;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01111111101010101010101010101010; //0 * NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b10000000000000000000000000000000; //inf * 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b10000000000000000000000000000000; //-inf * 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b01111111101010101010101010101010;	//inf * NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01111111101010101010101010101010; //-inf * NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b10000000000000000000000000000000; //NaN * 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b01111111100000000000000000000000;	//NaN * inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b11111111100000000000000000000000; //NaN * (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;


	///////////////////////////////////////////////////////
	////                    Divide                     ////
	///////////////////////////////////////////////////////
	op = 2'b11;
	//Normal cases
	inA=32'b01000010111010000000000000000000; inB=32'b01000000010000000000000000000000; //116 / 3
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01000010111010000000000000000000; inB=32'b11000000010000000000000000000000; //116 / (-3)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000010111010000000000000000000; inB=32'b01000000010000000000000000000000; //-116 / 3
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000010111010000000000000000000; inB=32'b11000000010000000000000000000000; //-116 / (-3)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b01000010111101101110100101111001; //0.69 / 123.456
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b11000010111101101110100101111001; //0.69 / (-123.456)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b01000010111101101110100101111001; //-0.69 / 123.456
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b11000010111101101110100101111001; //-0.69 / (-123.456)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b00111111001100001010001111010111; //0.69 / 0.69
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11000010111010000000000000000000; inB=32'b11000010111010000000000000000000; //-116 / (-116)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;

	//Zero cases
	inA=32'b00000000000000000000000000000000; inB=32'b01000000010000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01000000010000000000000000000000; // 0 / 3
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b11000000010000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b11000000010000000000000000000000; // 0 / (-3)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b10000000000000000000000000000000; // 0.69 / 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b10000000000000000000000000000000; // -0.69 / 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b10000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b10000000000000000000000000000000; // 0 / 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;

	//Infinity cases
	inA=32'b01111111100000000000000000000000; inB=32'b01000000010000000000000000000000;	// inf / 3
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01000000010000000000000000000000; // -inf / 3
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b11000000010000000000000000000000;	// inf / (-3)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b11000000010000000000000000000000; // -inf / (-3)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b01111111100000000000000000000000;	// 0.69 / inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b11111111100000000000000000000000; // 0.69 / (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b01111111100000000000000000000000;	// -0.69 / inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b11111111100000000000000000000000; // -0.69 / (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	// inf / inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b11111111100000000000000000000000;	// inf / (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	// -inf / inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b11111111100000000000000000000000; // -inf / (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;

	//Nan cases
	inA=32'b01111111101010101010101010101010; inB=32'b01000000010000000000000000000000;	// NaN / 3
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b11000000010000000000000000000000;	// NaN / (-3)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b01111111101010101010101010101010;	// 0.69 / NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b01111111101010101010101010101010;	// -0.69 / NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b01111111101010101010101010101010;	// NaN / NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;

	//Crossover
	inA=32'b00000000000000000000000000000000; inB=32'b01111111100000000000000000000000;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01111111100000000000000000000000; // 0 / inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b11111111100000000000000000000000;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b11111111100000000000000000000000; // 0 / (-inf)
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b01111111101010101010101010101010;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01111111101010101010101010101010; // 0 / NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b00000000000000000000000000000000;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b10000000000000000000000000000000; // inf / 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b00000000000000000000000000000000;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b10000000000000000000000000000000; // -inf / 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b01111111101010101010101010101010;	// inf / NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01111111101010101010101010101010; // -inf / NaN
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b00000000000000000000000000000000;	
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b10000000000000000000000000000000; // NaN / 0
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b01111111100000000000000000000000;	// NaN / inf
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b11111111100000000000000000000000; // NaN / (-inf)m
	#20 rst_n = 1 ; #260 ; rst_n = 0 ;
	$stop ;
end


always begin
	clk=~clk ;
	#10 ;
end

endmodule