module Mul24Bit(X,Y,Z);
input [23:0] X,Y;
output [47:0] Z;

//Hang Y0
assign Z[0]=X[0]&Y[0];

//Hang Y1
FullAdder fy1_0((X[1]&Y[0]),(X[0]&Y[1]),1'b0,Z[1],CY1_0);
FullAdder fy1_1((X[2]&Y[0]),(X[1]&Y[1]),CY1_0,Y1_0,CY1_1);
FullAdder fy1_2((X[3]&Y[0]),(X[2]&Y[1]),CY1_1,Y1_1,CY1_2);
FullAdder fy1_3((X[4]&Y[0]),(X[3]&Y[1]),CY1_2,Y1_2,CY1_3);
FullAdder fy1_4((X[5]&Y[0]),(X[4]&Y[1]),CY1_3,Y1_3,CY1_4);
FullAdder fy1_5((X[6]&Y[0]),(X[5]&Y[1]),CY1_4,Y1_4,CY1_5);
FullAdder fy1_6((X[7]&Y[0]),(X[6]&Y[1]),CY1_5,Y1_5,CY1_6);
FullAdder fy1_7((X[8]&Y[0]),(X[7]&Y[1]),CY1_6,Y1_6,CY1_7);
FullAdder fy1_8((X[9]&Y[0]),(X[8]&Y[1]),CY1_7,Y1_7,CY1_8);
FullAdder fy1_9((X[10]&Y[0]),(X[9]&Y[1]),CY1_8,Y1_8,CY1_9);
FullAdder fy1_10((X[11]&Y[0]),(X[10]&Y[1]),CY1_9,Y1_9,CY1_10);
FullAdder fy1_11((X[12]&Y[0]),(X[11]&Y[1]),CY1_10,Y1_10,CY1_11);
FullAdder fy1_12((X[13]&Y[0]),(X[12]&Y[1]),CY1_11,Y1_11,CY1_12);
FullAdder fy1_13((X[14]&Y[0]),(X[13]&Y[1]),CY1_12,Y1_12,CY1_13);
FullAdder fy1_14((X[15]&Y[0]),(X[14]&Y[1]),CY1_13,Y1_13,CY1_14);
FullAdder fy1_15((X[16]&Y[0]),(X[15]&Y[1]),CY1_14,Y1_14,CY1_15);
FullAdder fy1_16((X[17]&Y[0]),(X[16]&Y[1]),CY1_15,Y1_15,CY1_16);
FullAdder fy1_17((X[18]&Y[0]),(X[17]&Y[1]),CY1_16,Y1_16,CY1_17);
FullAdder fy1_18((X[19]&Y[0]),(X[18]&Y[1]),CY1_17,Y1_17,CY1_18);
FullAdder fy1_19((X[20]&Y[0]),(X[19]&Y[1]),CY1_18,Y1_18,CY1_19);
FullAdder fy1_20((X[21]&Y[0]),(X[20]&Y[1]),CY1_19,Y1_19,CY1_20);
FullAdder fy1_21((X[22]&Y[0]),(X[21]&Y[1]),CY1_20,Y1_20,CY1_21);
FullAdder fy1_22((X[23]&Y[0]),(X[22]&Y[1]),CY1_21,Y1_21,CY1_22);
FullAdder fy1_23(1'b0,(X[23]&Y[1]),CY1_22,Y1_22,Y2big);

//Hang Y2
FullAdder fy2_0(Y1_0,(X[0]&Y[2]),1'b0,Z[2],CY2_0);
FullAdder fy2_1(Y1_1,(X[1]&Y[2]),CY2_0,Y2_0,CY2_1);
FullAdder fy2_2(Y1_2,(X[2]&Y[2]),CY2_1,Y2_1,CY2_2);
FullAdder fy2_3(Y1_3,(X[3]&Y[2]),CY2_2,Y2_2,CY2_3);
FullAdder fy2_4(Y1_4,(X[4]&Y[2]),CY2_3,Y2_3,CY2_4);
FullAdder fy2_5(Y1_5,(X[5]&Y[2]),CY2_4,Y2_4,CY2_5);
FullAdder fy2_6(Y1_6,(X[6]&Y[2]),CY2_5,Y2_5,CY2_6);
FullAdder fy2_7(Y1_7,(X[7]&Y[2]),CY2_6,Y2_6,CY2_7);
FullAdder fy2_8(Y1_8,(X[8]&Y[2]),CY2_7,Y2_7,CY2_8);
FullAdder fy2_9(Y1_9,(X[9]&Y[2]),CY2_8,Y2_8,CY2_9);
FullAdder fy2_10(Y1_10,(X[10]&Y[2]),CY2_9,Y2_9,CY2_10);
FullAdder fy2_11(Y1_11,(X[11]&Y[2]),CY2_10,Y2_10,CY2_11);
FullAdder fy2_12(Y1_12,(X[12]&Y[2]),CY2_11,Y2_11,CY2_12);
FullAdder fy2_13(Y1_13,(X[13]&Y[2]),CY2_12,Y2_12,CY2_13);
FullAdder fy2_14(Y1_14,(X[14]&Y[2]),CY2_13,Y2_13,CY2_14);
FullAdder fy2_15(Y1_15,(X[15]&Y[2]),CY2_14,Y2_14,CY2_15);
FullAdder fy2_16(Y1_16,(X[16]&Y[2]),CY2_15,Y2_15,CY2_16);
FullAdder fy2_17(Y1_17,(X[17]&Y[2]),CY2_16,Y2_16,CY2_17);
FullAdder fy2_18(Y1_18,(X[18]&Y[2]),CY2_17,Y2_17,CY2_18);
FullAdder fy2_19(Y1_19,(X[19]&Y[2]),CY2_18,Y2_18,CY2_19);
FullAdder fy2_20(Y1_20,(X[20]&Y[2]),CY2_19,Y2_19,CY2_20);
FullAdder fy2_21(Y1_21,(X[21]&Y[2]),CY2_20,Y2_20,CY2_21);
FullAdder fy2_22(Y1_22,(X[22]&Y[2]),CY2_21,Y2_21,CY2_22);
FullAdder fy2_23(Y2big,(X[23]&Y[2]),CY2_22,Y2_22,Y3big);

//Hang Y3
FullAdder fy3_0(Y2_0,(X[0]&Y[3]),1'b0,Z[3],CY3_0);
FullAdder fy3_1(Y2_1,(X[1]&Y[3]),CY3_0,Y3_0,CY3_1);
FullAdder fy3_2(Y2_2,(X[2]&Y[3]),CY3_1,Y3_1,CY3_2);
FullAdder fy3_3(Y2_3,(X[3]&Y[3]),CY3_2,Y3_2,CY3_3);
FullAdder fy3_4(Y2_4,(X[4]&Y[3]),CY3_3,Y3_3,CY3_4);
FullAdder fy3_5(Y2_5,(X[5]&Y[3]),CY3_4,Y3_4,CY3_5);
FullAdder fy3_6(Y2_6,(X[6]&Y[3]),CY3_5,Y3_5,CY3_6);
FullAdder fy3_7(Y2_7,(X[7]&Y[3]),CY3_6,Y3_6,CY3_7);
FullAdder fy3_8(Y2_8,(X[8]&Y[3]),CY3_7,Y3_7,CY3_8);
FullAdder fy3_9(Y2_9,(X[9]&Y[3]),CY3_8,Y3_8,CY3_9);
FullAdder fy3_10(Y2_10,(X[10]&Y[3]),CY3_9,Y3_9,CY3_10);
FullAdder fy3_11(Y2_11,(X[11]&Y[3]),CY3_10,Y3_10,CY3_11);
FullAdder fy3_12(Y2_12,(X[12]&Y[3]),CY3_11,Y3_11,CY3_12);
FullAdder fy3_13(Y2_13,(X[13]&Y[3]),CY3_12,Y3_12,CY3_13);
FullAdder fy3_14(Y2_14,(X[14]&Y[3]),CY3_13,Y3_13,CY3_14);
FullAdder fy3_15(Y2_15,(X[15]&Y[3]),CY3_14,Y3_14,CY3_15);
FullAdder fy3_16(Y2_16,(X[16]&Y[3]),CY3_15,Y3_15,CY3_16);
FullAdder fy3_17(Y2_17,(X[17]&Y[3]),CY3_16,Y3_16,CY3_17);
FullAdder fy3_18(Y2_18,(X[18]&Y[3]),CY3_17,Y3_17,CY3_18);
FullAdder fy3_19(Y2_19,(X[19]&Y[3]),CY3_18,Y3_18,CY3_19);
FullAdder fy3_20(Y2_20,(X[20]&Y[3]),CY3_19,Y3_19,CY3_20);
FullAdder fy3_21(Y2_21,(X[21]&Y[3]),CY3_20,Y3_20,CY3_21);
FullAdder fy3_22(Y2_22,(X[22]&Y[3]),CY3_21,Y3_21,CY3_22);
FullAdder fy3_23(Y3big,(X[23]&Y[3]),CY3_22,Y3_22,Y4big);

//Hang Y4
FullAdder fy4_0(Y3_0,(X[0]&Y[4]),1'b0,Z[4],CY4_0);
FullAdder fy4_1(Y3_1,(X[1]&Y[4]),CY4_0,Y4_0,CY4_1);
FullAdder fy4_2(Y3_2,(X[2]&Y[4]),CY4_1,Y4_1,CY4_2);
FullAdder fy4_3(Y3_3,(X[3]&Y[4]),CY4_2,Y4_2,CY4_3);
FullAdder fy4_4(Y3_4,(X[4]&Y[4]),CY4_3,Y4_3,CY4_4);
FullAdder fy4_5(Y3_5,(X[5]&Y[4]),CY4_4,Y4_4,CY4_5);
FullAdder fy4_6(Y3_6,(X[6]&Y[4]),CY4_5,Y4_5,CY4_6);
FullAdder fy4_7(Y3_7,(X[7]&Y[4]),CY4_6,Y4_6,CY4_7);
FullAdder fy4_8(Y3_8,(X[8]&Y[4]),CY4_7,Y4_7,CY4_8);
FullAdder fy4_9(Y3_9,(X[9]&Y[4]),CY4_8,Y4_8,CY4_9);
FullAdder fy4_10(Y3_10,(X[10]&Y[4]),CY4_9,Y4_9,CY4_10);
FullAdder fy4_11(Y3_11,(X[11]&Y[4]),CY4_10,Y4_10,CY4_11);
FullAdder fy4_12(Y3_12,(X[12]&Y[4]),CY4_11,Y4_11,CY4_12);
FullAdder fy4_13(Y3_13,(X[13]&Y[4]),CY4_12,Y4_12,CY4_13);
FullAdder fy4_14(Y3_14,(X[14]&Y[4]),CY4_13,Y4_13,CY4_14);
FullAdder fy4_15(Y3_15,(X[15]&Y[4]),CY4_14,Y4_14,CY4_15);
FullAdder fy4_16(Y3_16,(X[16]&Y[4]),CY4_15,Y4_15,CY4_16);
FullAdder fy4_17(Y3_17,(X[17]&Y[4]),CY4_16,Y4_16,CY4_17);
FullAdder fy4_18(Y3_18,(X[18]&Y[4]),CY4_17,Y4_17,CY4_18);
FullAdder fy4_19(Y3_19,(X[19]&Y[4]),CY4_18,Y4_18,CY4_19);
FullAdder fy4_20(Y3_20,(X[20]&Y[4]),CY4_19,Y4_19,CY4_20);
FullAdder fy4_21(Y3_21,(X[21]&Y[4]),CY4_20,Y4_20,CY4_21);
FullAdder fy4_22(Y3_22,(X[22]&Y[4]),CY4_21,Y4_21,CY4_22);
FullAdder fy4_23(Y4big,(X[23]&Y[4]),CY4_22,Y4_22,Y5big);

//Hang Y5
FullAdder fy5_0(Y4_0,(X[0]&Y[5]),1'b0,Z[5],CY5_0);
FullAdder fy5_1(Y4_1,(X[1]&Y[5]),CY5_0,Y5_0,CY5_1);
FullAdder fy5_2(Y4_2,(X[2]&Y[5]),CY5_1,Y5_1,CY5_2);
FullAdder fy5_3(Y4_3,(X[3]&Y[5]),CY5_2,Y5_2,CY5_3);
FullAdder fy5_4(Y4_4,(X[4]&Y[5]),CY5_3,Y5_3,CY5_4);
FullAdder fy5_5(Y4_5,(X[5]&Y[5]),CY5_4,Y5_4,CY5_5);
FullAdder fy5_6(Y4_6,(X[6]&Y[5]),CY5_5,Y5_5,CY5_6);
FullAdder fy5_7(Y4_7,(X[7]&Y[5]),CY5_6,Y5_6,CY5_7);
FullAdder fy5_8(Y4_8,(X[8]&Y[5]),CY5_7,Y5_7,CY5_8);
FullAdder fy5_9(Y4_9,(X[9]&Y[5]),CY5_8,Y5_8,CY5_9);
FullAdder fy5_10(Y4_10,(X[10]&Y[5]),CY5_9,Y5_9,CY5_10);
FullAdder fy5_11(Y4_11,(X[11]&Y[5]),CY5_10,Y5_10,CY5_11);
FullAdder fy5_12(Y4_12,(X[12]&Y[5]),CY5_11,Y5_11,CY5_12);
FullAdder fy5_13(Y4_13,(X[13]&Y[5]),CY5_12,Y5_12,CY5_13);
FullAdder fy5_14(Y4_14,(X[14]&Y[5]),CY5_13,Y5_13,CY5_14);
FullAdder fy5_15(Y4_15,(X[15]&Y[5]),CY5_14,Y5_14,CY5_15);
FullAdder fy5_16(Y4_16,(X[16]&Y[5]),CY5_15,Y5_15,CY5_16);
FullAdder fy5_17(Y4_17,(X[17]&Y[5]),CY5_16,Y5_16,CY5_17);
FullAdder fy5_18(Y4_18,(X[18]&Y[5]),CY5_17,Y5_17,CY5_18);
FullAdder fy5_19(Y4_19,(X[19]&Y[5]),CY5_18,Y5_18,CY5_19);
FullAdder fy5_20(Y4_20,(X[20]&Y[5]),CY5_19,Y5_19,CY5_20);
FullAdder fy5_21(Y4_21,(X[21]&Y[5]),CY5_20,Y5_20,CY5_21);
FullAdder fy5_22(Y4_22,(X[22]&Y[5]),CY5_21,Y5_21,CY5_22);
FullAdder fy5_23(Y5big,(X[23]&Y[5]),CY5_22,Y5_22,Y6big);

//Hang Y6
FullAdder fy6_0(Y5_0,(X[0]&Y[6]),1'b0,Z[6],CY6_0);
FullAdder fy6_1(Y5_1,(X[1]&Y[6]),CY6_0,Y6_0,CY6_1);
FullAdder fy6_2(Y5_2,(X[2]&Y[6]),CY6_1,Y6_1,CY6_2);
FullAdder fy6_3(Y5_3,(X[3]&Y[6]),CY6_2,Y6_2,CY6_3);
FullAdder fy6_4(Y5_4,(X[4]&Y[6]),CY6_3,Y6_3,CY6_4);
FullAdder fy6_5(Y5_5,(X[5]&Y[6]),CY6_4,Y6_4,CY6_5);
FullAdder fy6_6(Y5_6,(X[6]&Y[6]),CY6_5,Y6_5,CY6_6);
FullAdder fy6_7(Y5_7,(X[7]&Y[6]),CY6_6,Y6_6,CY6_7);
FullAdder fy6_8(Y5_8,(X[8]&Y[6]),CY6_7,Y6_7,CY6_8);
FullAdder fy6_9(Y5_9,(X[9]&Y[6]),CY6_8,Y6_8,CY6_9);
FullAdder fy6_10(Y5_10,(X[10]&Y[6]),CY6_9,Y6_9,CY6_10);
FullAdder fy6_11(Y5_11,(X[11]&Y[6]),CY6_10,Y6_10,CY6_11);
FullAdder fy6_12(Y5_12,(X[12]&Y[6]),CY6_11,Y6_11,CY6_12);
FullAdder fy6_13(Y5_13,(X[13]&Y[6]),CY6_12,Y6_12,CY6_13);
FullAdder fy6_14(Y5_14,(X[14]&Y[6]),CY6_13,Y6_13,CY6_14);
FullAdder fy6_15(Y5_15,(X[15]&Y[6]),CY6_14,Y6_14,CY6_15);
FullAdder fy6_16(Y5_16,(X[16]&Y[6]),CY6_15,Y6_15,CY6_16);
FullAdder fy6_17(Y5_17,(X[17]&Y[6]),CY6_16,Y6_16,CY6_17);
FullAdder fy6_18(Y5_18,(X[18]&Y[6]),CY6_17,Y6_17,CY6_18);
FullAdder fy6_19(Y5_19,(X[19]&Y[6]),CY6_18,Y6_18,CY6_19);
FullAdder fy6_20(Y5_20,(X[20]&Y[6]),CY6_19,Y6_19,CY6_20);
FullAdder fy6_21(Y5_21,(X[21]&Y[6]),CY6_20,Y6_20,CY6_21);
FullAdder fy6_22(Y5_22,(X[22]&Y[6]),CY6_21,Y6_21,CY6_22);
FullAdder fy6_23(Y6big,(X[23]&Y[6]),CY6_22,Y6_22,Y7big);

//Hang Y7
FullAdder fy7_0(Y6_0,(X[0]&Y[7]),1'b0,Z[7],CY7_0);
FullAdder fy7_1(Y6_1,(X[1]&Y[7]),CY7_0,Y7_0,CY7_1);
FullAdder fy7_2(Y6_2,(X[2]&Y[7]),CY7_1,Y7_1,CY7_2);
FullAdder fy7_3(Y6_3,(X[3]&Y[7]),CY7_2,Y7_2,CY7_3);
FullAdder fy7_4(Y6_4,(X[4]&Y[7]),CY7_3,Y7_3,CY7_4);
FullAdder fy7_5(Y6_5,(X[5]&Y[7]),CY7_4,Y7_4,CY7_5);
FullAdder fy7_6(Y6_6,(X[6]&Y[7]),CY7_5,Y7_5,CY7_6);
FullAdder fy7_7(Y6_7,(X[7]&Y[7]),CY7_6,Y7_6,CY7_7);
FullAdder fy7_8(Y6_8,(X[8]&Y[7]),CY7_7,Y7_7,CY7_8);
FullAdder fy7_9(Y6_9,(X[9]&Y[7]),CY7_8,Y7_8,CY7_9);
FullAdder fy7_10(Y6_10,(X[10]&Y[7]),CY7_9,Y7_9,CY7_10);
FullAdder fy7_11(Y6_11,(X[11]&Y[7]),CY7_10,Y7_10,CY7_11);
FullAdder fy7_12(Y6_12,(X[12]&Y[7]),CY7_11,Y7_11,CY7_12);
FullAdder fy7_13(Y6_13,(X[13]&Y[7]),CY7_12,Y7_12,CY7_13);
FullAdder fy7_14(Y6_14,(X[14]&Y[7]),CY7_13,Y7_13,CY7_14);
FullAdder fy7_15(Y6_15,(X[15]&Y[7]),CY7_14,Y7_14,CY7_15);
FullAdder fy7_16(Y6_16,(X[16]&Y[7]),CY7_15,Y7_15,CY7_16);
FullAdder fy7_17(Y6_17,(X[17]&Y[7]),CY7_16,Y7_16,CY7_17);
FullAdder fy7_18(Y6_18,(X[18]&Y[7]),CY7_17,Y7_17,CY7_18);
FullAdder fy7_19(Y6_19,(X[19]&Y[7]),CY7_18,Y7_18,CY7_19);
FullAdder fy7_20(Y6_20,(X[20]&Y[7]),CY7_19,Y7_19,CY7_20);
FullAdder fy7_21(Y6_21,(X[21]&Y[7]),CY7_20,Y7_20,CY7_21);
FullAdder fy7_22(Y6_22,(X[22]&Y[7]),CY7_21,Y7_21,CY7_22);
FullAdder fy7_23(Y7big,(X[23]&Y[7]),CY7_22,Y7_22,Y8big);

//Hang Y8
FullAdder fy8_0(Y7_0,(X[0]&Y[8]),1'b0,Z[8],CY8_0);
FullAdder fy8_1(Y7_1,(X[1]&Y[8]),CY8_0,Y8_0,CY8_1);
FullAdder fy8_2(Y7_2,(X[2]&Y[8]),CY8_1,Y8_1,CY8_2);
FullAdder fy8_3(Y7_3,(X[3]&Y[8]),CY8_2,Y8_2,CY8_3);
FullAdder fy8_4(Y7_4,(X[4]&Y[8]),CY8_3,Y8_3,CY8_4);
FullAdder fy8_5(Y7_5,(X[5]&Y[8]),CY8_4,Y8_4,CY8_5);
FullAdder fy8_6(Y7_6,(X[6]&Y[8]),CY8_5,Y8_5,CY8_6);
FullAdder fy8_7(Y7_7,(X[7]&Y[8]),CY8_6,Y8_6,CY8_7);
FullAdder fy8_8(Y7_8,(X[8]&Y[8]),CY8_7,Y8_7,CY8_8);
FullAdder fy8_9(Y7_9,(X[9]&Y[8]),CY8_8,Y8_8,CY8_9);
FullAdder fy8_10(Y7_10,(X[10]&Y[8]),CY8_9,Y8_9,CY8_10);
FullAdder fy8_11(Y7_11,(X[11]&Y[8]),CY8_10,Y8_10,CY8_11);
FullAdder fy8_12(Y7_12,(X[12]&Y[8]),CY8_11,Y8_11,CY8_12);
FullAdder fy8_13(Y7_13,(X[13]&Y[8]),CY8_12,Y8_12,CY8_13);
FullAdder fy8_14(Y7_14,(X[14]&Y[8]),CY8_13,Y8_13,CY8_14);
FullAdder fy8_15(Y7_15,(X[15]&Y[8]),CY8_14,Y8_14,CY8_15);
FullAdder fy8_16(Y7_16,(X[16]&Y[8]),CY8_15,Y8_15,CY8_16);
FullAdder fy8_17(Y7_17,(X[17]&Y[8]),CY8_16,Y8_16,CY8_17);
FullAdder fy8_18(Y7_18,(X[18]&Y[8]),CY8_17,Y8_17,CY8_18);
FullAdder fy8_19(Y7_19,(X[19]&Y[8]),CY8_18,Y8_18,CY8_19);
FullAdder fy8_20(Y7_20,(X[20]&Y[8]),CY8_19,Y8_19,CY8_20);
FullAdder fy8_21(Y7_21,(X[21]&Y[8]),CY8_20,Y8_20,CY8_21);
FullAdder fy8_22(Y7_22,(X[22]&Y[8]),CY8_21,Y8_21,CY8_22);
FullAdder fy8_23(Y8big,(X[23]&Y[8]),CY8_22,Y8_22,Y9big);

//Hang Y9
FullAdder fy9_0(Y8_0,(X[0]&Y[9]),1'b0,Z[9],CY9_0);
FullAdder fy9_1(Y8_1,(X[1]&Y[9]),CY9_0,Y9_0,CY9_1);
FullAdder fy9_2(Y8_2,(X[2]&Y[9]),CY9_1,Y9_1,CY9_2);
FullAdder fy9_3(Y8_3,(X[3]&Y[9]),CY9_2,Y9_2,CY9_3);
FullAdder fy9_4(Y8_4,(X[4]&Y[9]),CY9_3,Y9_3,CY9_4);
FullAdder fy9_5(Y8_5,(X[5]&Y[9]),CY9_4,Y9_4,CY9_5);
FullAdder fy9_6(Y8_6,(X[6]&Y[9]),CY9_5,Y9_5,CY9_6);
FullAdder fy9_7(Y8_7,(X[7]&Y[9]),CY9_6,Y9_6,CY9_7);
FullAdder fy9_8(Y8_8,(X[8]&Y[9]),CY9_7,Y9_7,CY9_8);
FullAdder fy9_9(Y8_9,(X[9]&Y[9]),CY9_8,Y9_8,CY9_9);
FullAdder fy9_10(Y8_10,(X[10]&Y[9]),CY9_9,Y9_9,CY9_10);
FullAdder fy9_11(Y8_11,(X[11]&Y[9]),CY9_10,Y9_10,CY9_11);
FullAdder fy9_12(Y8_12,(X[12]&Y[9]),CY9_11,Y9_11,CY9_12);
FullAdder fy9_13(Y8_13,(X[13]&Y[9]),CY9_12,Y9_12,CY9_13);
FullAdder fy9_14(Y8_14,(X[14]&Y[9]),CY9_13,Y9_13,CY9_14);
FullAdder fy9_15(Y8_15,(X[15]&Y[9]),CY9_14,Y9_14,CY9_15);
FullAdder fy9_16(Y8_16,(X[16]&Y[9]),CY9_15,Y9_15,CY9_16);
FullAdder fy9_17(Y8_17,(X[17]&Y[9]),CY9_16,Y9_16,CY9_17);
FullAdder fy9_18(Y8_18,(X[18]&Y[9]),CY9_17,Y9_17,CY9_18);
FullAdder fy9_19(Y8_19,(X[19]&Y[9]),CY9_18,Y9_18,CY9_19);
FullAdder fy9_20(Y8_20,(X[20]&Y[9]),CY9_19,Y9_19,CY9_20);
FullAdder fy9_21(Y8_21,(X[21]&Y[9]),CY9_20,Y9_20,CY9_21);
FullAdder fy9_22(Y8_22,(X[22]&Y[9]),CY9_21,Y9_21,CY9_22);
FullAdder fy9_23(Y9big,(X[23]&Y[9]),CY9_22,Y9_22,Y10big);

//Hang Y10
FullAdder fy10_0(Y9_0,(X[0]&Y[10]),1'b0,Z[10],CY10_0);
FullAdder fy10_1(Y9_1,(X[1]&Y[10]),CY10_0,Y10_0,CY10_1);
FullAdder fy10_2(Y9_2,(X[2]&Y[10]),CY10_1,Y10_1,CY10_2);
FullAdder fy10_3(Y9_3,(X[3]&Y[10]),CY10_2,Y10_2,CY10_3);
FullAdder fy10_4(Y9_4,(X[4]&Y[10]),CY10_3,Y10_3,CY10_4);
FullAdder fy10_5(Y9_5,(X[5]&Y[10]),CY10_4,Y10_4,CY10_5);
FullAdder fy10_6(Y9_6,(X[6]&Y[10]),CY10_5,Y10_5,CY10_6);
FullAdder fy10_7(Y9_7,(X[7]&Y[10]),CY10_6,Y10_6,CY10_7);
FullAdder fy10_8(Y9_8,(X[8]&Y[10]),CY10_7,Y10_7,CY10_8);
FullAdder fy10_9(Y9_9,(X[9]&Y[10]),CY10_8,Y10_8,CY10_9);
FullAdder fy10_10(Y9_10,(X[10]&Y[10]),CY10_9,Y10_9,CY10_10);
FullAdder fy10_11(Y9_11,(X[11]&Y[10]),CY10_10,Y10_10,CY10_11);
FullAdder fy10_12(Y9_12,(X[12]&Y[10]),CY10_11,Y10_11,CY10_12);
FullAdder fy10_13(Y9_13,(X[13]&Y[10]),CY10_12,Y10_12,CY10_13);
FullAdder fy10_14(Y9_14,(X[14]&Y[10]),CY10_13,Y10_13,CY10_14);
FullAdder fy10_15(Y9_15,(X[15]&Y[10]),CY10_14,Y10_14,CY10_15);
FullAdder fy10_16(Y9_16,(X[16]&Y[10]),CY10_15,Y10_15,CY10_16);
FullAdder fy10_17(Y9_17,(X[17]&Y[10]),CY10_16,Y10_16,CY10_17);
FullAdder fy10_18(Y9_18,(X[18]&Y[10]),CY10_17,Y10_17,CY10_18);
FullAdder fy10_19(Y9_19,(X[19]&Y[10]),CY10_18,Y10_18,CY10_19);
FullAdder fy10_20(Y9_20,(X[20]&Y[10]),CY10_19,Y10_19,CY10_20);
FullAdder fy10_21(Y9_21,(X[21]&Y[10]),CY10_20,Y10_20,CY10_21);
FullAdder fy10_22(Y9_22,(X[22]&Y[10]),CY10_21,Y10_21,CY10_22);
FullAdder fy10_23(Y10big,(X[23]&Y[10]),CY10_22,Y10_22,Y11big);

//Hang Y11
FullAdder fy11_0(Y10_0,(X[0]&Y[11]),1'b0,Z[11],CY11_0);
FullAdder fy11_1(Y10_1,(X[1]&Y[11]),CY11_0,Y11_0,CY11_1);
FullAdder fy11_2(Y10_2,(X[2]&Y[11]),CY11_1,Y11_1,CY11_2);
FullAdder fy11_3(Y10_3,(X[3]&Y[11]),CY11_2,Y11_2,CY11_3);
FullAdder fy11_4(Y10_4,(X[4]&Y[11]),CY11_3,Y11_3,CY11_4);
FullAdder fy11_5(Y10_5,(X[5]&Y[11]),CY11_4,Y11_4,CY11_5);
FullAdder fy11_6(Y10_6,(X[6]&Y[11]),CY11_5,Y11_5,CY11_6);
FullAdder fy11_7(Y10_7,(X[7]&Y[11]),CY11_6,Y11_6,CY11_7);
FullAdder fy11_8(Y10_8,(X[8]&Y[11]),CY11_7,Y11_7,CY11_8);
FullAdder fy11_9(Y10_9,(X[9]&Y[11]),CY11_8,Y11_8,CY11_9);
FullAdder fy11_10(Y10_10,(X[10]&Y[11]),CY11_9,Y11_9,CY11_10);
FullAdder fy11_11(Y10_11,(X[11]&Y[11]),CY11_10,Y11_10,CY11_11);
FullAdder fy11_12(Y10_12,(X[12]&Y[11]),CY11_11,Y11_11,CY11_12);
FullAdder fy11_13(Y10_13,(X[13]&Y[11]),CY11_12,Y11_12,CY11_13);
FullAdder fy11_14(Y10_14,(X[14]&Y[11]),CY11_13,Y11_13,CY11_14);
FullAdder fy11_15(Y10_15,(X[15]&Y[11]),CY11_14,Y11_14,CY11_15);
FullAdder fy11_16(Y10_16,(X[16]&Y[11]),CY11_15,Y11_15,CY11_16);
FullAdder fy11_17(Y10_17,(X[17]&Y[11]),CY11_16,Y11_16,CY11_17);
FullAdder fy11_18(Y10_18,(X[18]&Y[11]),CY11_17,Y11_17,CY11_18);
FullAdder fy11_19(Y10_19,(X[19]&Y[11]),CY11_18,Y11_18,CY11_19);
FullAdder fy11_20(Y10_20,(X[20]&Y[11]),CY11_19,Y11_19,CY11_20);
FullAdder fy11_21(Y10_21,(X[21]&Y[11]),CY11_20,Y11_20,CY11_21);
FullAdder fy11_22(Y10_22,(X[22]&Y[11]),CY11_21,Y11_21,CY11_22);
FullAdder fy11_23(Y11big,(X[23]&Y[11]),CY11_22,Y11_22,Y12big);

//Hang Y12
FullAdder fy12_0(Y11_0,(X[0]&Y[12]),1'b0,Z[12],CY12_0);
FullAdder fy12_1(Y11_1,(X[1]&Y[12]),CY12_0,Y12_0,CY12_1);
FullAdder fy12_2(Y11_2,(X[2]&Y[12]),CY12_1,Y12_1,CY12_2);
FullAdder fy12_3(Y11_3,(X[3]&Y[12]),CY12_2,Y12_2,CY12_3);
FullAdder fy12_4(Y11_4,(X[4]&Y[12]),CY12_3,Y12_3,CY12_4);
FullAdder fy12_5(Y11_5,(X[5]&Y[12]),CY12_4,Y12_4,CY12_5);
FullAdder fy12_6(Y11_6,(X[6]&Y[12]),CY12_5,Y12_5,CY12_6);
FullAdder fy12_7(Y11_7,(X[7]&Y[12]),CY12_6,Y12_6,CY12_7);
FullAdder fy12_8(Y11_8,(X[8]&Y[12]),CY12_7,Y12_7,CY12_8);
FullAdder fy12_9(Y11_9,(X[9]&Y[12]),CY12_8,Y12_8,CY12_9);
FullAdder fy12_10(Y11_10,(X[10]&Y[12]),CY12_9,Y12_9,CY12_10);
FullAdder fy12_11(Y11_11,(X[11]&Y[12]),CY12_10,Y12_10,CY12_11);
FullAdder fy12_12(Y11_12,(X[12]&Y[12]),CY12_11,Y12_11,CY12_12);
FullAdder fy12_13(Y11_13,(X[13]&Y[12]),CY12_12,Y12_12,CY12_13);
FullAdder fy12_14(Y11_14,(X[14]&Y[12]),CY12_13,Y12_13,CY12_14);
FullAdder fy12_15(Y11_15,(X[15]&Y[12]),CY12_14,Y12_14,CY12_15);
FullAdder fy12_16(Y11_16,(X[16]&Y[12]),CY12_15,Y12_15,CY12_16);
FullAdder fy12_17(Y11_17,(X[17]&Y[12]),CY12_16,Y12_16,CY12_17);
FullAdder fy12_18(Y11_18,(X[18]&Y[12]),CY12_17,Y12_17,CY12_18);
FullAdder fy12_19(Y11_19,(X[19]&Y[12]),CY12_18,Y12_18,CY12_19);
FullAdder fy12_20(Y11_20,(X[20]&Y[12]),CY12_19,Y12_19,CY12_20);
FullAdder fy12_21(Y11_21,(X[21]&Y[12]),CY12_20,Y12_20,CY12_21);
FullAdder fy12_22(Y11_22,(X[22]&Y[12]),CY12_21,Y12_21,CY12_22);
FullAdder fy12_23(Y12big,(X[23]&Y[12]),CY12_22,Y12_22,Y13big);

//Hang Y13
FullAdder fy13_0(Y12_0,(X[0]&Y[13]),1'b0,Z[13],CY13_0);
FullAdder fy13_1(Y12_1,(X[1]&Y[13]),CY13_0,Y13_0,CY13_1);
FullAdder fy13_2(Y12_2,(X[2]&Y[13]),CY13_1,Y13_1,CY13_2);
FullAdder fy13_3(Y12_3,(X[3]&Y[13]),CY13_2,Y13_2,CY13_3);
FullAdder fy13_4(Y12_4,(X[4]&Y[13]),CY13_3,Y13_3,CY13_4);
FullAdder fy13_5(Y12_5,(X[5]&Y[13]),CY13_4,Y13_4,CY13_5);
FullAdder fy13_6(Y12_6,(X[6]&Y[13]),CY13_5,Y13_5,CY13_6);
FullAdder fy13_7(Y12_7,(X[7]&Y[13]),CY13_6,Y13_6,CY13_7);
FullAdder fy13_8(Y12_8,(X[8]&Y[13]),CY13_7,Y13_7,CY13_8);
FullAdder fy13_9(Y12_9,(X[9]&Y[13]),CY13_8,Y13_8,CY13_9);
FullAdder fy13_10(Y12_10,(X[10]&Y[13]),CY13_9,Y13_9,CY13_10);
FullAdder fy13_11(Y12_11,(X[11]&Y[13]),CY13_10,Y13_10,CY13_11);
FullAdder fy13_12(Y12_12,(X[12]&Y[13]),CY13_11,Y13_11,CY13_12);
FullAdder fy13_13(Y12_13,(X[13]&Y[13]),CY13_12,Y13_12,CY13_13);
FullAdder fy13_14(Y12_14,(X[14]&Y[13]),CY13_13,Y13_13,CY13_14);
FullAdder fy13_15(Y12_15,(X[15]&Y[13]),CY13_14,Y13_14,CY13_15);
FullAdder fy13_16(Y12_16,(X[16]&Y[13]),CY13_15,Y13_15,CY13_16);
FullAdder fy13_17(Y12_17,(X[17]&Y[13]),CY13_16,Y13_16,CY13_17);
FullAdder fy13_18(Y12_18,(X[18]&Y[13]),CY13_17,Y13_17,CY13_18);
FullAdder fy13_19(Y12_19,(X[19]&Y[13]),CY13_18,Y13_18,CY13_19);
FullAdder fy13_20(Y12_20,(X[20]&Y[13]),CY13_19,Y13_19,CY13_20);
FullAdder fy13_21(Y12_21,(X[21]&Y[13]),CY13_20,Y13_20,CY13_21);
FullAdder fy13_22(Y12_22,(X[22]&Y[13]),CY13_21,Y13_21,CY13_22);
FullAdder fy13_23(Y13big,(X[23]&Y[13]),CY13_22,Y13_22,Y14big);

//Hang Y14
FullAdder fy14_0(Y13_0,(X[0]&Y[14]),1'b0,Z[14],CY14_0);
FullAdder fy14_1(Y13_1,(X[1]&Y[14]),CY14_0,Y14_0,CY14_1);
FullAdder fy14_2(Y13_2,(X[2]&Y[14]),CY14_1,Y14_1,CY14_2);
FullAdder fy14_3(Y13_3,(X[3]&Y[14]),CY14_2,Y14_2,CY14_3);
FullAdder fy14_4(Y13_4,(X[4]&Y[14]),CY14_3,Y14_3,CY14_4);
FullAdder fy14_5(Y13_5,(X[5]&Y[14]),CY14_4,Y14_4,CY14_5);
FullAdder fy14_6(Y13_6,(X[6]&Y[14]),CY14_5,Y14_5,CY14_6);
FullAdder fy14_7(Y13_7,(X[7]&Y[14]),CY14_6,Y14_6,CY14_7);
FullAdder fy14_8(Y13_8,(X[8]&Y[14]),CY14_7,Y14_7,CY14_8);
FullAdder fy14_9(Y13_9,(X[9]&Y[14]),CY14_8,Y14_8,CY14_9);
FullAdder fy14_10(Y13_10,(X[10]&Y[14]),CY14_9,Y14_9,CY14_10);
FullAdder fy14_11(Y13_11,(X[11]&Y[14]),CY14_10,Y14_10,CY14_11);
FullAdder fy14_12(Y13_12,(X[12]&Y[14]),CY14_11,Y14_11,CY14_12);
FullAdder fy14_13(Y13_13,(X[13]&Y[14]),CY14_12,Y14_12,CY14_13);
FullAdder fy14_14(Y13_14,(X[14]&Y[14]),CY14_13,Y14_13,CY14_14);
FullAdder fy14_15(Y13_15,(X[15]&Y[14]),CY14_14,Y14_14,CY14_15);
FullAdder fy14_16(Y13_16,(X[16]&Y[14]),CY14_15,Y14_15,CY14_16);
FullAdder fy14_17(Y13_17,(X[17]&Y[14]),CY14_16,Y14_16,CY14_17);
FullAdder fy14_18(Y13_18,(X[18]&Y[14]),CY14_17,Y14_17,CY14_18);
FullAdder fy14_19(Y13_19,(X[19]&Y[14]),CY14_18,Y14_18,CY14_19);
FullAdder fy14_20(Y13_20,(X[20]&Y[14]),CY14_19,Y14_19,CY14_20);
FullAdder fy14_21(Y13_21,(X[21]&Y[14]),CY14_20,Y14_20,CY14_21);
FullAdder fy14_22(Y13_22,(X[22]&Y[14]),CY14_21,Y14_21,CY14_22);
FullAdder fy14_23(Y14big,(X[23]&Y[14]),CY14_22,Y14_22,Y15big);

//Hang Y15
FullAdder fy15_0(Y14_0,(X[0]&Y[15]),1'b0,Z[15],CY15_0);
FullAdder fy15_1(Y14_1,(X[1]&Y[15]),CY15_0,Y15_0,CY15_1);
FullAdder fy15_2(Y14_2,(X[2]&Y[15]),CY15_1,Y15_1,CY15_2);
FullAdder fy15_3(Y14_3,(X[3]&Y[15]),CY15_2,Y15_2,CY15_3);
FullAdder fy15_4(Y14_4,(X[4]&Y[15]),CY15_3,Y15_3,CY15_4);
FullAdder fy15_5(Y14_5,(X[5]&Y[15]),CY15_4,Y15_4,CY15_5);
FullAdder fy15_6(Y14_6,(X[6]&Y[15]),CY15_5,Y15_5,CY15_6);
FullAdder fy15_7(Y14_7,(X[7]&Y[15]),CY15_6,Y15_6,CY15_7);
FullAdder fy15_8(Y14_8,(X[8]&Y[15]),CY15_7,Y15_7,CY15_8);
FullAdder fy15_9(Y14_9,(X[9]&Y[15]),CY15_8,Y15_8,CY15_9);
FullAdder fy15_10(Y14_10,(X[10]&Y[15]),CY15_9,Y15_9,CY15_10);
FullAdder fy15_11(Y14_11,(X[11]&Y[15]),CY15_10,Y15_10,CY15_11);
FullAdder fy15_12(Y14_12,(X[12]&Y[15]),CY15_11,Y15_11,CY15_12);
FullAdder fy15_13(Y14_13,(X[13]&Y[15]),CY15_12,Y15_12,CY15_13);
FullAdder fy15_14(Y14_14,(X[14]&Y[15]),CY15_13,Y15_13,CY15_14);
FullAdder fy15_15(Y14_15,(X[15]&Y[15]),CY15_14,Y15_14,CY15_15);
FullAdder fy15_16(Y14_16,(X[16]&Y[15]),CY15_15,Y15_15,CY15_16);
FullAdder fy15_17(Y14_17,(X[17]&Y[15]),CY15_16,Y15_16,CY15_17);
FullAdder fy15_18(Y14_18,(X[18]&Y[15]),CY15_17,Y15_17,CY15_18);
FullAdder fy15_19(Y14_19,(X[19]&Y[15]),CY15_18,Y15_18,CY15_19);
FullAdder fy15_20(Y14_20,(X[20]&Y[15]),CY15_19,Y15_19,CY15_20);
FullAdder fy15_21(Y14_21,(X[21]&Y[15]),CY15_20,Y15_20,CY15_21);
FullAdder fy15_22(Y14_22,(X[22]&Y[15]),CY15_21,Y15_21,CY15_22);
FullAdder fy15_23(Y15big,(X[23]&Y[15]),CY15_22,Y15_22,Y16big);

//Hang Y16
FullAdder fy16_0(Y15_0,(X[0]&Y[16]),1'b0,Z[16],CY16_0);
FullAdder fy16_1(Y15_1,(X[1]&Y[16]),CY16_0,Y16_0,CY16_1);
FullAdder fy16_2(Y15_2,(X[2]&Y[16]),CY16_1,Y16_1,CY16_2);
FullAdder fy16_3(Y15_3,(X[3]&Y[16]),CY16_2,Y16_2,CY16_3);
FullAdder fy16_4(Y15_4,(X[4]&Y[16]),CY16_3,Y16_3,CY16_4);
FullAdder fy16_5(Y15_5,(X[5]&Y[16]),CY16_4,Y16_4,CY16_5);
FullAdder fy16_6(Y15_6,(X[6]&Y[16]),CY16_5,Y16_5,CY16_6);
FullAdder fy16_7(Y15_7,(X[7]&Y[16]),CY16_6,Y16_6,CY16_7);
FullAdder fy16_8(Y15_8,(X[8]&Y[16]),CY16_7,Y16_7,CY16_8);
FullAdder fy16_9(Y15_9,(X[9]&Y[16]),CY16_8,Y16_8,CY16_9);
FullAdder fy16_10(Y15_10,(X[10]&Y[16]),CY16_9,Y16_9,CY16_10);
FullAdder fy16_11(Y15_11,(X[11]&Y[16]),CY16_10,Y16_10,CY16_11);
FullAdder fy16_12(Y15_12,(X[12]&Y[16]),CY16_11,Y16_11,CY16_12);
FullAdder fy16_13(Y15_13,(X[13]&Y[16]),CY16_12,Y16_12,CY16_13);
FullAdder fy16_14(Y15_14,(X[14]&Y[16]),CY16_13,Y16_13,CY16_14);
FullAdder fy16_15(Y15_15,(X[15]&Y[16]),CY16_14,Y16_14,CY16_15);
FullAdder fy16_16(Y15_16,(X[16]&Y[16]),CY16_15,Y16_15,CY16_16);
FullAdder fy16_17(Y15_17,(X[17]&Y[16]),CY16_16,Y16_16,CY16_17);
FullAdder fy16_18(Y15_18,(X[18]&Y[16]),CY16_17,Y16_17,CY16_18);
FullAdder fy16_19(Y15_19,(X[19]&Y[16]),CY16_18,Y16_18,CY16_19);
FullAdder fy16_20(Y15_20,(X[20]&Y[16]),CY16_19,Y16_19,CY16_20);
FullAdder fy16_21(Y15_21,(X[21]&Y[16]),CY16_20,Y16_20,CY16_21);
FullAdder fy16_22(Y15_22,(X[22]&Y[16]),CY16_21,Y16_21,CY16_22);
FullAdder fy16_23(Y16big,(X[23]&Y[16]),CY16_22,Y16_22,Y17big);

//Hang Y17
FullAdder fy17_0(Y16_0,(X[0]&Y[17]),1'b0,Z[17],CY17_0);
FullAdder fy17_1(Y16_1,(X[1]&Y[17]),CY17_0,Y17_0,CY17_1);
FullAdder fy17_2(Y16_2,(X[2]&Y[17]),CY17_1,Y17_1,CY17_2);
FullAdder fy17_3(Y16_3,(X[3]&Y[17]),CY17_2,Y17_2,CY17_3);
FullAdder fy17_4(Y16_4,(X[4]&Y[17]),CY17_3,Y17_3,CY17_4);
FullAdder fy17_5(Y16_5,(X[5]&Y[17]),CY17_4,Y17_4,CY17_5);
FullAdder fy17_6(Y16_6,(X[6]&Y[17]),CY17_5,Y17_5,CY17_6);
FullAdder fy17_7(Y16_7,(X[7]&Y[17]),CY17_6,Y17_6,CY17_7);
FullAdder fy17_8(Y16_8,(X[8]&Y[17]),CY17_7,Y17_7,CY17_8);
FullAdder fy17_9(Y16_9,(X[9]&Y[17]),CY17_8,Y17_8,CY17_9);
FullAdder fy17_10(Y16_10,(X[10]&Y[17]),CY17_9,Y17_9,CY17_10);
FullAdder fy17_11(Y16_11,(X[11]&Y[17]),CY17_10,Y17_10,CY17_11);
FullAdder fy17_12(Y16_12,(X[12]&Y[17]),CY17_11,Y17_11,CY17_12);
FullAdder fy17_13(Y16_13,(X[13]&Y[17]),CY17_12,Y17_12,CY17_13);
FullAdder fy17_14(Y16_14,(X[14]&Y[17]),CY17_13,Y17_13,CY17_14);
FullAdder fy17_15(Y16_15,(X[15]&Y[17]),CY17_14,Y17_14,CY17_15);
FullAdder fy17_16(Y16_16,(X[16]&Y[17]),CY17_15,Y17_15,CY17_16);
FullAdder fy17_17(Y16_17,(X[17]&Y[17]),CY17_16,Y17_16,CY17_17);
FullAdder fy17_18(Y16_18,(X[18]&Y[17]),CY17_17,Y17_17,CY17_18);
FullAdder fy17_19(Y16_19,(X[19]&Y[17]),CY17_18,Y17_18,CY17_19);
FullAdder fy17_20(Y16_20,(X[20]&Y[17]),CY17_19,Y17_19,CY17_20);
FullAdder fy17_21(Y16_21,(X[21]&Y[17]),CY17_20,Y17_20,CY17_21);
FullAdder fy17_22(Y16_22,(X[22]&Y[17]),CY17_21,Y17_21,CY17_22);
FullAdder fy17_23(Y17big,(X[23]&Y[17]),CY17_22,Y17_22,Y18big);

//Hang Y18
FullAdder fy18_0(Y17_0,(X[0]&Y[18]),1'b0,Z[18],CY18_0);
FullAdder fy18_1(Y17_1,(X[1]&Y[18]),CY18_0,Y18_0,CY18_1);
FullAdder fy18_2(Y17_2,(X[2]&Y[18]),CY18_1,Y18_1,CY18_2);
FullAdder fy18_3(Y17_3,(X[3]&Y[18]),CY18_2,Y18_2,CY18_3);
FullAdder fy18_4(Y17_4,(X[4]&Y[18]),CY18_3,Y18_3,CY18_4);
FullAdder fy18_5(Y17_5,(X[5]&Y[18]),CY18_4,Y18_4,CY18_5);
FullAdder fy18_6(Y17_6,(X[6]&Y[18]),CY18_5,Y18_5,CY18_6);
FullAdder fy18_7(Y17_7,(X[7]&Y[18]),CY18_6,Y18_6,CY18_7);
FullAdder fy18_8(Y17_8,(X[8]&Y[18]),CY18_7,Y18_7,CY18_8);
FullAdder fy18_9(Y17_9,(X[9]&Y[18]),CY18_8,Y18_8,CY18_9);
FullAdder fy18_10(Y17_10,(X[10]&Y[18]),CY18_9,Y18_9,CY18_10);
FullAdder fy18_11(Y17_11,(X[11]&Y[18]),CY18_10,Y18_10,CY18_11);
FullAdder fy18_12(Y17_12,(X[12]&Y[18]),CY18_11,Y18_11,CY18_12);
FullAdder fy18_13(Y17_13,(X[13]&Y[18]),CY18_12,Y18_12,CY18_13);
FullAdder fy18_14(Y17_14,(X[14]&Y[18]),CY18_13,Y18_13,CY18_14);
FullAdder fy18_15(Y17_15,(X[15]&Y[18]),CY18_14,Y18_14,CY18_15);
FullAdder fy18_16(Y17_16,(X[16]&Y[18]),CY18_15,Y18_15,CY18_16);
FullAdder fy18_17(Y17_17,(X[17]&Y[18]),CY18_16,Y18_16,CY18_17);
FullAdder fy18_18(Y17_18,(X[18]&Y[18]),CY18_17,Y18_17,CY18_18);
FullAdder fy18_19(Y17_19,(X[19]&Y[18]),CY18_18,Y18_18,CY18_19);
FullAdder fy18_20(Y17_20,(X[20]&Y[18]),CY18_19,Y18_19,CY18_20);
FullAdder fy18_21(Y17_21,(X[21]&Y[18]),CY18_20,Y18_20,CY18_21);
FullAdder fy18_22(Y17_22,(X[22]&Y[18]),CY18_21,Y18_21,CY18_22);
FullAdder fy18_23(Y18big,(X[23]&Y[18]),CY18_22,Y18_22,Y19big);

//Hang Y19
FullAdder fy19_0(Y18_0,(X[0]&Y[19]),1'b0,Z[19],CY19_0);
FullAdder fy19_1(Y18_1,(X[1]&Y[19]),CY19_0,Y19_0,CY19_1);
FullAdder fy19_2(Y18_2,(X[2]&Y[19]),CY19_1,Y19_1,CY19_2);
FullAdder fy19_3(Y18_3,(X[3]&Y[19]),CY19_2,Y19_2,CY19_3);
FullAdder fy19_4(Y18_4,(X[4]&Y[19]),CY19_3,Y19_3,CY19_4);
FullAdder fy19_5(Y18_5,(X[5]&Y[19]),CY19_4,Y19_4,CY19_5);
FullAdder fy19_6(Y18_6,(X[6]&Y[19]),CY19_5,Y19_5,CY19_6);
FullAdder fy19_7(Y18_7,(X[7]&Y[19]),CY19_6,Y19_6,CY19_7);
FullAdder fy19_8(Y18_8,(X[8]&Y[19]),CY19_7,Y19_7,CY19_8);
FullAdder fy19_9(Y18_9,(X[9]&Y[19]),CY19_8,Y19_8,CY19_9);
FullAdder fy19_10(Y18_10,(X[10]&Y[19]),CY19_9,Y19_9,CY19_10);
FullAdder fy19_11(Y18_11,(X[11]&Y[19]),CY19_10,Y19_10,CY19_11);
FullAdder fy19_12(Y18_12,(X[12]&Y[19]),CY19_11,Y19_11,CY19_12);
FullAdder fy19_13(Y18_13,(X[13]&Y[19]),CY19_12,Y19_12,CY19_13);
FullAdder fy19_14(Y18_14,(X[14]&Y[19]),CY19_13,Y19_13,CY19_14);
FullAdder fy19_15(Y18_15,(X[15]&Y[19]),CY19_14,Y19_14,CY19_15);
FullAdder fy19_16(Y18_16,(X[16]&Y[19]),CY19_15,Y19_15,CY19_16);
FullAdder fy19_17(Y18_17,(X[17]&Y[19]),CY19_16,Y19_16,CY19_17);
FullAdder fy19_18(Y18_18,(X[18]&Y[19]),CY19_17,Y19_17,CY19_18);
FullAdder fy19_19(Y18_19,(X[19]&Y[19]),CY19_18,Y19_18,CY19_19);
FullAdder fy19_20(Y18_20,(X[20]&Y[19]),CY19_19,Y19_19,CY19_20);
FullAdder fy19_21(Y18_21,(X[21]&Y[19]),CY19_20,Y19_20,CY19_21);
FullAdder fy19_22(Y18_22,(X[22]&Y[19]),CY19_21,Y19_21,CY19_22);
FullAdder fy19_23(Y19big,(X[23]&Y[19]),CY19_22,Y19_22,Y20big);

//Hang Y20
FullAdder fy20_0(Y19_0,(X[0]&Y[20]),1'b0,Z[20],CY20_0);
FullAdder fy20_1(Y19_1,(X[1]&Y[20]),CY20_0,Y20_0,CY20_1);
FullAdder fy20_2(Y19_2,(X[2]&Y[20]),CY20_1,Y20_1,CY20_2);
FullAdder fy20_3(Y19_3,(X[3]&Y[20]),CY20_2,Y20_2,CY20_3);
FullAdder fy20_4(Y19_4,(X[4]&Y[20]),CY20_3,Y20_3,CY20_4);
FullAdder fy20_5(Y19_5,(X[5]&Y[20]),CY20_4,Y20_4,CY20_5);
FullAdder fy20_6(Y19_6,(X[6]&Y[20]),CY20_5,Y20_5,CY20_6);
FullAdder fy20_7(Y19_7,(X[7]&Y[20]),CY20_6,Y20_6,CY20_7);
FullAdder fy20_8(Y19_8,(X[8]&Y[20]),CY20_7,Y20_7,CY20_8);
FullAdder fy20_9(Y19_9,(X[9]&Y[20]),CY20_8,Y20_8,CY20_9);
FullAdder fy20_10(Y19_10,(X[10]&Y[20]),CY20_9,Y20_9,CY20_10);
FullAdder fy20_11(Y19_11,(X[11]&Y[20]),CY20_10,Y20_10,CY20_11);
FullAdder fy20_12(Y19_12,(X[12]&Y[20]),CY20_11,Y20_11,CY20_12);
FullAdder fy20_13(Y19_13,(X[13]&Y[20]),CY20_12,Y20_12,CY20_13);
FullAdder fy20_14(Y19_14,(X[14]&Y[20]),CY20_13,Y20_13,CY20_14);
FullAdder fy20_15(Y19_15,(X[15]&Y[20]),CY20_14,Y20_14,CY20_15);
FullAdder fy20_16(Y19_16,(X[16]&Y[20]),CY20_15,Y20_15,CY20_16);
FullAdder fy20_17(Y19_17,(X[17]&Y[20]),CY20_16,Y20_16,CY20_17);
FullAdder fy20_18(Y19_18,(X[18]&Y[20]),CY20_17,Y20_17,CY20_18);
FullAdder fy20_19(Y19_19,(X[19]&Y[20]),CY20_18,Y20_18,CY20_19);
FullAdder fy20_20(Y19_20,(X[20]&Y[20]),CY20_19,Y20_19,CY20_20);
FullAdder fy20_21(Y19_21,(X[21]&Y[20]),CY20_20,Y20_20,CY20_21);
FullAdder fy20_22(Y19_22,(X[22]&Y[20]),CY20_21,Y20_21,CY20_22);
FullAdder fy20_23(Y20big,(X[23]&Y[20]),CY20_22,Y20_22,Y21big);

//Hang Y21
FullAdder fy21_0(Y20_0,(X[0]&Y[21]),1'b0,Z[21],CY21_0);
FullAdder fy21_1(Y20_1,(X[1]&Y[21]),CY21_0,Y21_0,CY21_1);
FullAdder fy21_2(Y20_2,(X[2]&Y[21]),CY21_1,Y21_1,CY21_2);
FullAdder fy21_3(Y20_3,(X[3]&Y[21]),CY21_2,Y21_2,CY21_3);
FullAdder fy21_4(Y20_4,(X[4]&Y[21]),CY21_3,Y21_3,CY21_4);
FullAdder fy21_5(Y20_5,(X[5]&Y[21]),CY21_4,Y21_4,CY21_5);
FullAdder fy21_6(Y20_6,(X[6]&Y[21]),CY21_5,Y21_5,CY21_6);
FullAdder fy21_7(Y20_7,(X[7]&Y[21]),CY21_6,Y21_6,CY21_7);
FullAdder fy21_8(Y20_8,(X[8]&Y[21]),CY21_7,Y21_7,CY21_8);
FullAdder fy21_9(Y20_9,(X[9]&Y[21]),CY21_8,Y21_8,CY21_9);
FullAdder fy21_10(Y20_10,(X[10]&Y[21]),CY21_9,Y21_9,CY21_10);
FullAdder fy21_11(Y20_11,(X[11]&Y[21]),CY21_10,Y21_10,CY21_11);
FullAdder fy21_12(Y20_12,(X[12]&Y[21]),CY21_11,Y21_11,CY21_12);
FullAdder fy21_13(Y20_13,(X[13]&Y[21]),CY21_12,Y21_12,CY21_13);
FullAdder fy21_14(Y20_14,(X[14]&Y[21]),CY21_13,Y21_13,CY21_14);
FullAdder fy21_15(Y20_15,(X[15]&Y[21]),CY21_14,Y21_14,CY21_15);
FullAdder fy21_16(Y20_16,(X[16]&Y[21]),CY21_15,Y21_15,CY21_16);
FullAdder fy21_17(Y20_17,(X[17]&Y[21]),CY21_16,Y21_16,CY21_17);
FullAdder fy21_18(Y20_18,(X[18]&Y[21]),CY21_17,Y21_17,CY21_18);
FullAdder fy21_19(Y20_19,(X[19]&Y[21]),CY21_18,Y21_18,CY21_19);
FullAdder fy21_20(Y20_20,(X[20]&Y[21]),CY21_19,Y21_19,CY21_20);
FullAdder fy21_21(Y20_21,(X[21]&Y[21]),CY21_20,Y21_20,CY21_21);
FullAdder fy21_22(Y20_22,(X[22]&Y[21]),CY21_21,Y21_21,CY21_22);
FullAdder fy21_23(Y21big,(X[23]&Y[21]),CY21_22,Y21_22,Y22big);

//Hang Y22
FullAdder fy22_0(Y21_0,(X[0]&Y[22]),1'b0,Z[22],CY22_0);
FullAdder fy22_1(Y21_1,(X[1]&Y[22]),CY22_0,Y22_0,CY22_1);
FullAdder fy22_2(Y21_2,(X[2]&Y[22]),CY22_1,Y22_1,CY22_2);
FullAdder fy22_3(Y21_3,(X[3]&Y[22]),CY22_2,Y22_2,CY22_3);
FullAdder fy22_4(Y21_4,(X[4]&Y[22]),CY22_3,Y22_3,CY22_4);
FullAdder fy22_5(Y21_5,(X[5]&Y[22]),CY22_4,Y22_4,CY22_5);
FullAdder fy22_6(Y21_6,(X[6]&Y[22]),CY22_5,Y22_5,CY22_6);
FullAdder fy22_7(Y21_7,(X[7]&Y[22]),CY22_6,Y22_6,CY22_7);
FullAdder fy22_8(Y21_8,(X[8]&Y[22]),CY22_7,Y22_7,CY22_8);
FullAdder fy22_9(Y21_9,(X[9]&Y[22]),CY22_8,Y22_8,CY22_9);
FullAdder fy22_10(Y21_10,(X[10]&Y[22]),CY22_9,Y22_9,CY22_10);
FullAdder fy22_11(Y21_11,(X[11]&Y[22]),CY22_10,Y22_10,CY22_11);
FullAdder fy22_12(Y21_12,(X[12]&Y[22]),CY22_11,Y22_11,CY22_12);
FullAdder fy22_13(Y21_13,(X[13]&Y[22]),CY22_12,Y22_12,CY22_13);
FullAdder fy22_14(Y21_14,(X[14]&Y[22]),CY22_13,Y22_13,CY22_14);
FullAdder fy22_15(Y21_15,(X[15]&Y[22]),CY22_14,Y22_14,CY22_15);
FullAdder fy22_16(Y21_16,(X[16]&Y[22]),CY22_15,Y22_15,CY22_16);
FullAdder fy22_17(Y21_17,(X[17]&Y[22]),CY22_16,Y22_16,CY22_17);
FullAdder fy22_18(Y21_18,(X[18]&Y[22]),CY22_17,Y22_17,CY22_18);
FullAdder fy22_19(Y21_19,(X[19]&Y[22]),CY22_18,Y22_18,CY22_19);
FullAdder fy22_20(Y21_20,(X[20]&Y[22]),CY22_19,Y22_19,CY22_20);
FullAdder fy22_21(Y21_21,(X[21]&Y[22]),CY22_20,Y22_20,CY22_21);
FullAdder fy22_22(Y21_22,(X[22]&Y[22]),CY22_21,Y22_21,CY22_22);
FullAdder fy22_23(Y22big,(X[23]&Y[22]),CY22_22,Y22_22,Y23big);

//Hang Y23
FullAdder fy23_0(Y22_0,(X[0]&Y[23]),1'b0,Z[23],CY23_0);
FullAdder fy23_1(Y22_1,(X[1]&Y[23]),CY23_0,Z[24],CY23_1);
FullAdder fy23_2(Y22_2,(X[2]&Y[23]),CY23_1,Z[25],CY23_2);
FullAdder fy23_3(Y22_3,(X[3]&Y[23]),CY23_2,Z[26],CY23_3);
FullAdder fy23_4(Y22_4,(X[4]&Y[23]),CY23_3,Z[27],CY23_4);
FullAdder fy23_5(Y22_5,(X[5]&Y[23]),CY23_4,Z[28],CY23_5);
FullAdder fy23_6(Y22_6,(X[6]&Y[23]),CY23_5,Z[29],CY23_6);
FullAdder fy23_7(Y22_7,(X[7]&Y[23]),CY23_6,Z[30],CY23_7);
FullAdder fy23_8(Y22_8,(X[8]&Y[23]),CY23_7,Z[31],CY23_8);
FullAdder fy23_9(Y22_9,(X[9]&Y[23]),CY23_8,Z[32],CY23_9);
FullAdder fy23_10(Y22_10,(X[10]&Y[23]),CY23_9,Z[33],CY23_10);
FullAdder fy23_11(Y22_11,(X[11]&Y[23]),CY23_10,Z[34],CY23_11);
FullAdder fy23_12(Y22_12,(X[12]&Y[23]),CY23_11,Z[35],CY23_12);
FullAdder fy23_13(Y22_13,(X[13]&Y[23]),CY23_12,Z[36],CY23_13);
FullAdder fy23_14(Y22_14,(X[14]&Y[23]),CY23_13,Z[37],CY23_14);
FullAdder fy23_15(Y22_15,(X[15]&Y[23]),CY23_14,Z[38],CY23_15);
FullAdder fy23_16(Y22_16,(X[16]&Y[23]),CY23_15,Z[39],CY23_16);
FullAdder fy23_17(Y22_17,(X[17]&Y[23]),CY23_16,Z[40],CY23_17);
FullAdder fy23_18(Y22_18,(X[18]&Y[23]),CY23_17,Z[41],CY23_18);
FullAdder fy23_19(Y22_19,(X[19]&Y[23]),CY23_18,Z[42],CY23_19);
FullAdder fy23_20(Y22_20,(X[20]&Y[23]),CY23_19,Z[43],CY23_20);
FullAdder fy23_21(Y22_21,(X[21]&Y[23]),CY23_20,Z[44],CY23_21);
FullAdder fy23_22(Y22_22,(X[22]&Y[23]),CY23_21,Z[45],CY23_22);
FullAdder fy23_23(Y23big,(X[23]&Y[23]),CY23_22,Z[46],Z[47]);


endmodule


