module fa (
	output	s, c,
	input		x, y, z
);
wire		w;

assign	w = x ^ y ;
assign	s = w ^ z ;
assign	c = (w & z) | (x & y) ;

endmodule
//====================================

module csa_26b (x,y,z,s,cout);
	output [25:0] 	s;
	output cout;
	input  [25:0]	x, y, z;

wire	[25:0]	s1, c1 ;
wire	[24:0]	w ;

fa		pre_00	(s1[00], c1[00], x[00], y[00], z[00]) ;
fa		pre_01	(s1[01], c1[01], x[01], y[01], z[01]) ;
fa		pre_02	(s1[02], c1[02], x[02], y[02], z[02]) ;
fa		pre_03	(s1[03], c1[03], x[03], y[03], z[03]) ;
fa		pre_04	(s1[04], c1[04], x[04], y[04], z[04]) ;
fa		pre_05	(s1[05], c1[05], x[05], y[05], z[05]) ;
fa		pre_06	(s1[06], c1[06], x[06], y[06], z[06]) ;
fa		pre_07	(s1[07], c1[07], x[07], y[07], z[07]) ;
fa		pre_08	(s1[08], c1[08], x[08], y[08], z[08]) ;
fa		pre_09	(s1[09], c1[09], x[09], y[09], z[09]) ;
fa		pre_10	(s1[10], c1[10], x[10], y[10], z[10]) ;
fa		pre_11	(s1[11], c1[11], x[11], y[11], z[11]) ;
fa		pre_12	(s1[12], c1[12], x[12], y[12], z[12]) ;
fa		pre_13	(s1[13], c1[13], x[13], y[13], z[13]) ;
fa		pre_14	(s1[14], c1[14], x[14], y[14], z[14]) ;
fa		pre_15	(s1[15], c1[15], x[15], y[15], z[15]) ;
fa		pre_16	(s1[16], c1[16], x[16], y[16], z[16]) ;
fa		pre_17	(s1[17], c1[17], x[17], y[17], z[17]) ;
fa		pre_18	(s1[18], c1[18], x[18], y[18], z[18]) ;
fa		pre_19	(s1[19], c1[19], x[19], y[19], z[19]) ;
fa		pre_20	(s1[20], c1[20], x[20], y[20], z[20]) ;
fa		pre_21	(s1[21], c1[21], x[21], y[21], z[21]) ;
fa		pre_22	(s1[22], c1[22], x[22], y[22], z[22]) ;
fa		pre_23	(s1[23], c1[23], x[23], y[23], z[23]) ;
fa		pre_24	(s1[24], c1[24], x[24], y[24], z[24]) ;
fa		pre_25	(s1[25], c1[25], x[25], y[25], z[25]) ;

assign		s[00] = s1[00] ;
assign		cout 	= w[24] ;
fa		b_01		(s[01], w[00], s1[01], c1[00], 1'b0) ;
fa		b_02		(s[02], w[01], s1[02], c1[01], w[00]) ;
fa		b_03		(s[03], w[02], s1[03], c1[02], w[01]) ;
fa		b_04		(s[04], w[03], s1[04], c1[03], w[02]) ;
fa		b_05		(s[05], w[04], s1[05], c1[04], w[03]) ;
fa		b_06		(s[06], w[05], s1[06], c1[05], w[04]) ;
fa		b_07		(s[07], w[06], s1[07], c1[06], w[05]) ;
fa		b_08		(s[08], w[07], s1[08], c1[07], w[06]) ;
fa		b_09		(s[09], w[08], s1[09], c1[08], w[07]) ;
fa		b_10		(s[10], w[09], s1[10], c1[09], w[08]) ;
fa		b_11		(s[11], w[10], s1[11], c1[10], w[09]) ;
fa		b_12		(s[12], w[11], s1[12], c1[11], w[10]) ;
fa		b_13		(s[13], w[12], s1[13], c1[12], w[11]) ;
fa		b_14		(s[14], w[13], s1[14], c1[13], w[12]) ;
fa		b_15		(s[15], w[14], s1[15], c1[14], w[13]) ;
fa		b_16		(s[16], w[15], s1[16], c1[15], w[14]) ;
fa		b_17		(s[17], w[16], s1[17], c1[16], w[15]) ;
fa		b_18		(s[18], w[17], s1[18], c1[17], w[16]) ;
fa		b_19		(s[19], w[18], s1[19], c1[18], w[17]) ;
fa		b_20		(s[20], w[19], s1[20], c1[19], w[18]) ;
fa		b_21		(s[21], w[20], s1[21], c1[20], w[19]) ;
fa		b_22		(s[22], w[21], s1[22], c1[21], w[20]) ;
fa		b_23		(s[23], w[22], s1[23], c1[22], w[21]) ;
fa		b_24		(s[24], w[23], s1[24], c1[23], w[22]) ;
fa		b_25		(s[25], w[24], s1[25], c1[24], w[23]) ;

endmodule
