module Multiplication_tb;
reg [31:0] inA, inB;
reg clk;
wire [31:0] out;

Multiplication M_tb(inA,inB,clk,out);
always begin #10 clk=~clk; end

initial begin 
//Normal cases
#0 clk=1;inA=32'b00111111110000000000000000000000; inB=32'b01000010101110010101110000101001; //1.5 * 92.68
#20 inA=32'b00111111110000000000000000000000; inB=32'b11000010101110010101110000101001; //1.5 * (-92.68)
#20 inA=32'b10111111110000000000000000000000; inB=32'b01000010101110010101110000101001; //-1.5 * 92.68
#20 inA=32'b10111111110000000000000000000000; inB=32'b11000010101110010101110000101001; //-1.5 * (-92.68)
//Zero cases
#20 inA=32'b00000000000000000000000000000000; inB=32'b01000010101110010101110000101001; 
#20 inA=32'b10000000000000000000000000000000; inB=32'b01000010101110010101110000101001; //0 * 92.68
#20 inA=32'b00000000000000000000000000000000; inB=32'b11000010101110010101110000101001; 
#20 inA=32'b10000000000000000000000000000000; inB=32'b11000010101110010101110000101001; //0 * (-92.68)
#20 inA=32'b00111111110000000000000000000000; inB=32'b00000000000000000000000000000000;
#20 inA=32'b00111111110000000000000000000000; inB=32'b10000000000000000000000000000000; //1.5 * 0
#20 inA=32'b10111111110000000000000000000000; inB=32'b00000000000000000000000000000000;
#20 inA=32'b10111111110000000000000000000000; inB=32'b10000000000000000000000000000000; //-1.5 * 0
#20 inA=32'b00000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
#20 inA=32'b00000000000000000000000000000000; inB=32'b10000000000000000000000000000000;
#20 inA=32'b10000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
#20 inA=32'b10000000000000000000000000000000; inB=32'b10000000000000000000000000000000; //0 * 0
//Infinity cases
#20 inA=32'b01111111100000000000000000000000; inB=32'b01000010101110010101110000101001; //inf * 92.68
#20 inA=32'b11111111100000000000000000000000; inB=32'b01000010101110010101110000101001; //-inf * 92.68
#20 inA=32'b01111111100000000000000000000000; inB=32'b11000010101110010101110000101001; //inf * (-92.68)
#20 inA=32'b11111111100000000000000000000000; inB=32'b11000010101110010101110000101001; //-inf * (-92.68)
#20 inA=32'b00111111110000000000000000000000; inB=32'b01111111100000000000000000000000; //1.5 * inf
#20 inA=32'b00111111110000000000000000000000; inB=32'b11111111100000000000000000000000; //1.5 * (-inf)
#20 inA=32'b10111111110000000000000000000000; inB=32'b01111111100000000000000000000000; //-1.5 * inf
#20 inA=32'b10111111110000000000000000000000; inB=32'b11111111100000000000000000000000; //-1.5 * (-inf)
#20 inA=32'b01111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	//inf * inf
#20 inA=32'b01111111100000000000000000000000; inB=32'b11111111100000000000000000000000;	//inf * (-inf)
#20 inA=32'b11111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	//-inf * inf
#20 inA=32'b11111111100000000000000000000000; inB=32'b11111111100000000000000000000000;	//-inf * (-inf)
//NaN cases
#20 inA=32'b00111111110000000000000000000000; inB=32'b01111111101010101010101010101010; //1.5 * NaN
#20 inA=32'b10111111110000000000000000000000; inB=32'b01111111101010101010101010101010; //-1.5 * NaN
#20 inA=32'b01111111101010101010101010101010; inB=32'b01000010101110010101110000101001; //NaN * 92.68
#20 inA=32'b01111111101010101010101010101010; inB=32'b11000010101110010101110000101001; //NaN * (-92.68)
#20 inA=32'b01111111101010101010101010101010; inB=32'b01111111101010101010101010101010; //NaN * NaN
//Crossover cases
#20 inA=32'b00000000000000000000000000000000; inB=32'b01111111100000000000000000000000;
#20 inA=32'b10000000000000000000000000000000; inB=32'b01111111100000000000000000000000; //0 * inf
#20 inA=32'b00000000000000000000000000000000; inB=32'b11111111100000000000000000000000;
#20 inA=32'b10000000000000000000000000000000; inB=32'b11111111100000000000000000000000; //0 * (-inf)
#20 inA=32'b00000000000000000000000000000000; inB=32'b01111111101010101010101010101010;
#20 inA=32'b10000000000000000000000000000000; inB=32'b01111111101010101010101010101010; //0 * NaN
#20 inA=32'b01111111100000000000000000000000; inB=32'b00000000000000000000000000000000;
#20 inA=32'b01111111100000000000000000000000; inB=32'b10000000000000000000000000000000; //inf * 0
#20 inA=32'b11111111100000000000000000000000; inB=32'b00000000000000000000000000000000;
#20 inA=32'b11111111100000000000000000000000; inB=32'b10000000000000000000000000000000; //-inf * 0
#20 inA=32'b01111111100000000000000000000000; inB=32'b01111111101010101010101010101010;	//inf * NaN
#20 inA=32'b11111111100000000000000000000000; inB=32'b01111111101010101010101010101010; //-inf * NaN
#20 inA=32'b01111111101010101010101010101010; inB=32'b00000000000000000000000000000000;
#20 inA=32'b01111111101010101010101010101010; inB=32'b10000000000000000000000000000000; //NaN * 0
#20 inA=32'b01111111101010101010101010101010; inB=32'b01111111100000000000000000000000;	//NaN * inf
#20 inA=32'b01111111101010101010101010101010; inB=32'b11111111100000000000000000000000; //NaN * (-inf)
#20; $stop;
end

endmodule	