module AddSub_tb;

reg [31:0] inA,inB;
reg op;
wire [31:0] out;

AddSub AS0(inA,inB,op,out);

initial begin
//Test for normal numbers

#20 inA=32'b01000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//7.5 + 1.46
#20 inA=32'b01000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//7.5 + (-1.46)
#20 inA=32'b01000000111100000000000000000000;inB=32'b11000001000101110101110000101001; op=0;	//7.5 + (-9.46)
#20 inA=32'b11000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//(-7.5)+1.46
#20 inA=32'b11000000111100000000000000000000;inB=32'b01000001000101110101110000101001; op=0;	//(-7.5)+9.46
#20 inA=32'b11000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//(-7.5)+(-1.46)
#20 inA=32'b01000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//7.5 - 1.46
#20 inA=32'b01000000111100000000000000000000;inB=32'b01000001000101110101110000101001; op=1;	//7.5 - 9.46
#20 inA=32'b01000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//7.5 - (-1.46)
#20 inA=32'b11000000111100000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//(-7.5)-1.46
#20 inA=32'b11000000111100000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//-7.5 - (-1.46)
#20 inA=32'b11000000111100000000000000000000;inB=32'b11000001000101110101110000101001; op=1;	//-7.5 - (-9.46)
#20 inA=32'b01000000111100000000000000000000;inB=32'b01000000111100000000000000000000; op=1;	//7.5 - 7.5
#20 inA=32'b01000000111100000000000000000000;inB=32'b11000000111100000000000000000000; op=0;	//7.5 + (-7.5)
#20 inA=32'b11000000111100000000000000000000;inB=32'b01000000111100000000000000000000; op=0;	//-7.5 + 7.5
#20 inA=32'b11000000111100000000000000000000;inB=32'b11000000111100000000000000000000; op=1;	//-7.5 - (-7.5)

//Test for zero
#20 inA=32'b01000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
#20 inA=32'b01000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=0; 	//7.5+0
#20 inA=32'b01000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
#20 inA=32'b01000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=1; 	//7.5-0
#20 inA=32'b11000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
#20 inA=32'b11000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=0; 	//-7.5+0
#20 inA=32'b11000000111100000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
#20 inA=32'b11000000111100000000000000000000;inB=32'b10000000000000000000000000000000; op=1; 	//-7.5-0
#20 inA=32'b00000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;
#20 inA=32'b10000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//0+1.46
#20 inA=32'b00000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;
#20 inA=32'b10000000000000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//0-1.46
#20 inA=32'b00000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;
#20 inA=32'b10000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//0+(-1.46)
#20 inA=32'b00000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;
#20 inA=32'b10000000000000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//0-(-1.46)
#20 inA=32'b00000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
#20 inA=32'b00000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;
#20 inA=32'b10000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
#20 inA=32'b10000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;	//0+0
#20 inA=32'b00000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
#20 inA=32'b00000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;
#20 inA=32'b10000000000000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
#20 inA=32'b10000000000000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;	//0-0

//Test for infinity
#20 inA=32'b01000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//7.5+inf
#20 inA=32'b01000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//7.5-inf
#20 inA=32'b01000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//7.5+(-inf)
#20 inA=32'b01000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//7.5-(-inf)
#20 inA=32'b11000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//-7.5+inf
#20 inA=32'b11000000111100000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//-7.5-inf
#20 inA=32'b11000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//-7.5+(-inf)
#20 inA=32'b11000000111100000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//-7.5-(-inf)
#20 inA=32'b01111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//inf+1.46
#20 inA=32'b01111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//inf-1.46
#20 inA=32'b01111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//inf+(-1.46)
#20 inA=32'b01111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//inf-(-1.46)
#20 inA=32'b11111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=0;	//-inf+1.46
#20 inA=32'b11111111100000000000000000000000;inB=32'b00111111101110101110000101001000; op=1;	//-inf-1.46
#20 inA=32'b11111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=0;	//-inf+(-1.46)
#20 inA=32'b11111111100000000000000000000000;inB=32'b10111111101110101110000101001000; op=1;	//-inf-(-1.46)
#20 inA=32'b01111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//inf+inf
#20 inA=32'b01111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//inf-inf
#20 inA=32'b01111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//inf+(-inf)
#20 inA=32'b01111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//inf-(-inf)
#20 inA=32'b11111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//-inf+inf
#20 inA=32'b11111111100000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//-inf-inf
#20 inA=32'b11111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//-inf+(-inf)
#20 inA=32'b11111111100000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//-inf-(-inf)

//Test for NaN
#20 inA=32'b01000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//7.5+NaN
#20 inA=32'b01000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//7.5+NaN
#20 inA=32'b11000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//-7.5+NaN
#20 inA=32'b11000000111100000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//-7.5-NaN
#20 inA=32'b01111111101010101010101010101010;inB=32'b00111111101110101110000101001000; op=0;	//NaN+1.46
#20 inA=32'b01111111101010101010101010101010;inB=32'b00111111101110101110000101001000; op=1;	//NaN-1.46
#20 inA=32'b01111111101010101010101010101010;inB=32'b10111111101110101110000101001000; op=0;	//NaN+(-1.46)
#20 inA=32'b01111111101010101010101010101010;inB=32'b10111111101110101110000101001000; op=1;	//NaN-(-1.46)
#20 inA=32'b01111111101010101010101010101010;inB=32'b01111111101010101010101010101010; op=0;	//NaN+NaN
#20 inA=32'b01111111101010101010101010101010;inB=32'b01111111101010101010101010101010; op=1;	//NaN-NaN

//Crossover: Nan and inf and zero
#20 inA=32'b00000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;
#20 inA=32'b10000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=0;	//0+inf
#20 inA=32'b00000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;
#20 inA=32'b10000000000000000000000000000000;inB=32'b01111111100000000000000000000000; op=1;	//0+inf
#20 inA=32'b00000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;
#20 inA=32'b10000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=0;	//0+(-inf)
#20 inA=32'b00000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;
#20 inA=32'b10000000000000000000000000000000;inB=32'b11111111100000000000000000000000; op=1;	//0-(-inf)
#20 inA=32'b01111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
#20 inA=32'b01111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;	//inf+0
#20 inA=32'b01111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
#20 inA=32'b01111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;	//inf-0
#20 inA=32'b11111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=0;
#20 inA=32'b11111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=0;	//-inf+0
#20 inA=32'b11111111100000000000000000000000;inB=32'b00000000000000000000000000000000; op=1;
#20 inA=32'b11111111100000000000000000000000;inB=32'b10000000000000000000000000000000; op=1;	//-inf-0
#20 inA=32'b00000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	
#20 inA=32'b10000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//0+NaN
#20 inA=32'b00000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	
#20 inA=32'b10000000000000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//0-NaN
#20 inA=32'b01111111101010101010101010101010;inB=32'b00000000000000000000000000000000; op=0;	
#20 inA=32'b01111111101010101010101010101010;inB=32'b10000000000000000000000000000000; op=0;	//NaN+0
#20 inA=32'b01111111101010101010101010101010;inB=32'b00000000000000000000000000000000; op=1;	
#20 inA=32'b01111111101010101010101010101010;inB=32'b10000000000000000000000000000000; op=1;	//NaN-0
#20 inA=32'b01111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//inf+NaN
#20 inA=32'b01111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//inf-NaN
#20 inA=32'b11111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=0;	//-inf+NaN
#20 inA=32'b11111111100000000000000000000000;inB=32'b01111111101010101010101010101010; op=1;	//-inf-NaN
#20 inA=32'b01111111101010101010101010101010;inB=32'b01111111100000000000000000000000; op=0;	//NaN+inf
#20 inA=32'b01111111101010101010101010101010;inB=32'b01111111100000000000000000000000; op=1;	//NaN-inf
#20 inA=32'b01111111101010101010101010101010;inB=32'b11111111100000000000000000000000; op=0;	//NaN+(-inf)
#20 inA=32'b01111111101010101010101010101010;inB=32'b11111111100000000000000000000000; op=1;	//NaN-(-inf)

#20; $stop;

end

endmodule