module slct_q (mul_n3, mul_n2, mul_n1, mul_0, mul_1, mul_2, mul_3, finish, s, d, clk, n_rst, en);

output			mul_n3, mul_n2, mul_n1, mul_0, mul_1, mul_2, mul_3, finish ;
input			clk, n_rst, en ;
input	[4:0]	s, d ;

//assign mul_n3 =   (s[4] &&  s[3] &&  s[2] && !s[1] && !s[0] &&  d[3] &&  d[2])                  ||
// 		     		(s[4] &&  s[3] &&  s[2] && !s[1] &&           d[3] &&  d[2] &&  d[1])         ||
// 		     		(s[4] &&  s[3] && !s[2] &&  s[1] && !s[0] &&  d[3] &&           d[1])         ||
// 		     		(s[4] &&  s[3] && !s[2] &&  s[1] &&           d[3] &&  d[2])                  ||
// 		     		(s[4] &&  s[3] && !s[2] &&  s[1] &&           d[3] &&           d[1] && d[0]) ||
// 		     		(s[4] &&  s[3] && !s[2] && !s[1] &&  s[0] &&  d[3] &&          !d[1] && d[0]) ||
// 		     		(s[4] &&  s[3] && !s[2] && !s[1] && !s[0] &&  d[3] && !d[2])                  ||
// 		     		(s[4] &&  s[3] && !s[2] && !s[1] &&           d[3] && !d[2] &&  d[1])         ||
// 		     		(s[4] &&  s[3] && !s[2] &&           s[0] &&  d[3] &&  d[2] && !d[1])         ||
// 		     		(s[4] &&  s[3] &&           s[1] && !s[0] &&  d[3] &&  d[2] &&  d[1])         ||
// 		     		(s[4] &&  s[3] &&           s[1] &&           d[3] &&  d[2] &&  d[1] && d[0]) ||
// 		     		(s[4] &&  s[3] &&          !s[1] &&  s[0] &&  d[3] &&  d[2] && !d[1] && d[0]) ||
// 		     		(s[4] && !s[3] &&  s[2] &&  s[1] &&  s[0] &&  d[3] && !d[2] && !d[1]) ;

// updated
assign mul_n3 = (s[4]  &&  s[3]  &&  s[2]  && !s[1]  && !s[0]  &&  d[3]  &&  d[2])                     ||
				(s[4]  &&  s[3]  &&  s[2]  && !s[1]  &&            d[3]  &&  d[2]  &&  d[1])           ||
				(s[4]  &&  s[3]  && !s[2]  &&  s[1]  && !s[0]  &&  d[3]  &&            d[1])           ||
				(s[4]  &&  s[3]  && !s[2]  &&  s[1]  &&            d[3]  &&  d[2])                     ||
				(s[4]  &&  s[3]  && !s[2]  &&  s[1]  &&            d[3]  &&            d[1]  &&  d[0]) ||
				(s[4]  &&  s[3]  && !s[2]  && !s[1]  &&  s[0]  &&  d[3]  &&           !d[1]  &&  d[0]) ||
				(s[4]  &&  s[3]  && !s[2]  && !s[1]  && !s[0]  &&  d[3]  && !d[2])                     ||
				(s[4]  &&  s[3]  && !s[2]  && !s[1]  &&            d[3]  && !d[2]  &&  d[1])           ||
				(s[4]  &&  s[3]  && !s[2]  &&            s[0]  &&  d[3]  &&  d[2]  && !d[1])           ||
				(s[4]  &&  s[3]  &&            s[1]  && !s[0]  &&  d[3]  &&  d[2]  &&  d[1])           ||
				(s[4]  &&  s[3]  &&            s[1]  &&            d[3]  &&  d[2]  &&  d[1]  &&  d[0]) ||
				(s[4]  &&  s[3]  &&           !s[1]  &&  s[0]  &&  d[3]  &&  d[2]  && !d[1]  &&  d[0]) ||
				(s[4]  && !s[3]  &&  s[2]  &&  s[1]  &&  s[0]  &&  d[3]  && !d[2]  && !d[1])           ||
				(s[4]  && !s[3]  &&  s[2]  &&  s[1]  &&            d[3]  && !d[2]  && !d[1]  && !d[0]) ;


//
// assign mul_n2 = 
// 				(s[4] &&  s[3] && !s[2] && !s[1] && !s[0] &&  d[3] &&  d[2])                  ||
// 				(s[4] &&  s[3] && !s[2] && !s[1] &&           d[3] &&  d[2] &&  d[1])         ||
// 				(s[4] && !s[3] &&  s[2] &&  s[1] &&  s[0] &&  d[3] &&           d[1])         ||
// 				(s[4] && !s[3] &&  s[2] &&  s[1] &&           d[3] &&  d[2] && !d[1])         ||
// 				(s[4] && !s[3] &&  s[2] &&  s[1] &&           d[3] && !d[2] &&  d[1])         ||
// 				(s[4] && !s[3] &&  s[2] && !s[1] &&  s[0] &&  d[3] && !d[2])                  ||
// 				(s[4] && !s[3] &&  s[2] &&          !s[0] &&  d[3] && !d[2] && !d[1]) ;
// updated
assign mul_n2 = 
				(s[4]  &&  s[3]  && !s[2]  && !s[1]  && !s[0]  &&  d[3]  &&  d[2])                    ||
				(s[4]  &&  s[3]  && !s[2]  && !s[1]  &&            d[3]  &&  d[2]  &&  d[1])          ||
				(s[4]  && !s[3]  &&  s[2]  &&  s[1]  &&  s[0]  &&  d[3]  &&            d[1])          ||
				(s[4]  && !s[3]  &&  s[2]  &&  s[1]  &&            d[3]  &&  d[2]  && !d[1])          ||
				(s[4]  && !s[3]  &&  s[2]  &&  s[1]  &&            d[3]  && !d[2]  &&  d[1])          ||
				(s[4]  && !s[3]  &&  s[2]  && !s[1]  &&            d[3]  && !d[2]  && !d[1])          ||
				(s[4]  && !s[3]  &&  s[2]  &&            s[0]  &&  d[3]  && !d[2]  &&  d[1])          ||
				(s[4]  && !s[3]  &&  s[2]  &&           !s[0]  &&  d[3]  && !d[2]  && !d[1]  &&  d[0]) ;

assign mul_n1 = 
				(s[4] && !s[3] &&  s[2] && !s[1] && !s[0] &&  d[3] &&           d[1])         ||
				(s[4] && !s[3] &&  s[2] && !s[1] &&           d[3] &&   d[2])                 ||
				(s[4] && !s[3] &&  s[2] &&          !s[0] &&  d[3] &&   d[2] && d[1])         ||
				(s[4] && !s[3] && !s[2] &&  s[1] &&  s[0] &&  d[3])                           ||
				(s[4] && !s[3] && !s[2] &&  s[1] &&           d[3] &&  !d[2]) ;

assign mul_0  = 
				(s[4] && !s[3] && !s[2] && !s[1] &&           d[3])                           ||
				(s[4] && !s[3] && !s[2] &&          !s[0] &&  d[3] &&  d[2])                  ||
				(        !s[3] && !s[2] && !s[1] && !s[0] &&  d[3])                           ||
				(        !s[3] && !s[2] && !s[1] &&           d[3] &&  d[2] &&  d[1])         ||
				(        !s[3] && !s[2] && !s[1] &&           d[3] &&  d[2] &&         d[0]) ;

assign mul_1  = 
				( !s[4] && !s[3] &&  s[2] && !s[1] && !s[0] &&  d[3] &&  d[2] &&  d[1])          ||
				( !s[4] && !s[3] &&  s[2] && !s[1] && !s[0] &&  d[3] &&  d[2] &&           d[0]) ||
				( !s[4] && !s[3] &&  s[2] && !s[1] &&           d[3] &&  d[2] &&  d[1] &&  d[0]) ||
				( !s[4] && !s[3] && !s[2] &&  s[1] && !s[0] &&  d[3] )                           ||
				( !s[4] && !s[3] && !s[2] &&  s[1] &&           d[3] &&  d[2])                   ||
				( !s[4] && !s[3] && !s[2] &&  s[1] &&           d[3] &&           d[1] &&  d[0]) ||
				( !s[4] && !s[3] && !s[2] && !s[1] &&  s[0] &&  d[3] && !d[2])                   ||
				( !s[4] && !s[3] && !s[2] && !s[1] &&  s[0] &&  d[3] &&          !d[1] && !d[0]) ;

// assign mul_2  = 
// 				( !s[4] &&  s[3] && !s[2] && !s[1] && !s[0] &&  d[3] &&  d[2] &&  d[1] &&  d[0])    ||
// 				( !s[4] && !s[3] &&  s[2] &&  s[1] &&           d[3] &&  d[2] &&  d[1])             ||
// 				( !s[4] && !s[3] &&  s[2] &&  s[1]          &&  d[3] &&  d[2] &&           d[0])    ||
// 				( !s[4] && !s[3] &&  s[2] && !s[1] &&  s[0] &&  d[3] &&                   !d[0])    ||
// 				( !s[4] && !s[3] &&  s[2] && !s[1] &&           d[3] && !d[2] )                     ||
// 				( !s[4] && !s[3] &&  s[2] &&           s[0] &&  d[3] &&  d[2] && !d[1] &&  d[0])    ||
// 				( !s[4] && !s[3] &&  s[2] &&          !s[0] &&  d[3] &&  d[2] && !d[1] && !d[0])    ||
// 				( !s[4] && !s[3] &&  s[2] &&          !s[0] &&  d[3] && !d[2] &&  d[1] &&  d[0])    ||
// 				( !s[4] && !s[3] && !s[2] &&  s[1] &&  s[0] &&  d[3] && !d[2] && !d[1])             ||
// 				( !s[4] && !s[3] && !s[2] &&  s[1] &&  s[0] &&  d[3] && !d[2] &&          !d[0]) ;

// updated
assign mul_2 = 
				( !s[4]  &&  s[3]  && !s[2]  && !s[1]  && !s[0]  &&  d[3] &&  d[2] &&  d[1] &&  d[0])||
				( !s[4]  && !s[3]  &&  s[2]  &&  s[1]  && !s[0]  &&  d[3] &&  d[2])                  ||
				( !s[4]  && !s[3]  &&  s[2]  &&  s[1]  && !s[0]  &&  d[3] &&           d[1] &&  d[0])||
				( !s[4]  && !s[3]  &&  s[2]  &&  s[1]  &&            d[3] &&  d[2] &&  d[1])         ||
				( !s[4]  && !s[3]  &&  s[2]  && !s[1]  && !s[0]  &&  d[3] && !d[2])                  ||
				( !s[4]  && !s[3]  &&  s[2]  && !s[1]  &&            d[3] &&  d[2] && !d[1] && !d[0])||
				( !s[4]  && !s[3]  &&  s[2]  && !s[1]  &&            d[3] && !d[2] &&  d[1])         ||
				( !s[4]  && !s[3]  &&  s[2]  &&            s[0]  &&  d[3] &&  d[2] &&  d[1] && !d[0])||
				( !s[4]  && !s[3]  &&  s[2]  &&            s[0]  &&  d[3] &&  d[2] && !d[1] &&  d[0])||
				( !s[4]  && !s[3]  && !s[2]  &&  s[1]  &&  s[0]  &&  d[3] && !d[2] && !d[1])         ||
				( !s[4]  && !s[3]  && !s[2]  &&  s[1]  &&  s[0]  &&  d[3] && !d[2] &&          !d[0]) ;

// assign mul_3  = 
// 				( !s[4] &&  s[3] &&  s[2] &&          !s[0] &&  d[3] &&  d[2] &&  d[1])            ||
// 				( !s[4] &&  s[3] && !s[2] &&  s[1] && !s[0] &&  d[3] && !d[2] && !d[1] && !d[0])   ||
// 				( !s[4] &&  s[3] && !s[2] &&  s[1] &&           d[3] &&  d[2] )                    ||
// 				( !s[4] &&  s[3] && !s[2] && !s[1] &&  s[0] &&  d[3] &&           d[1])            ||
// 				( !s[4] &&  s[3] && !s[2] && !s[1] && !s[0] &&  d[3] &&                   !d[0])   ||
// 				( !s[4] &&  s[3] && !s[2] && !s[1] &&           d[3] &&          !d[1] &&  d[0])   ||
// 				( !s[4] &&  s[3] && !s[2] &&           s[0] &&  d[3] &&  d[2] )                    ||
// 				( !s[4] &&  s[3] && !s[2] &&                    d[3] && !d[2] &&  d[1] &&  d[0])   ||
// 				( !s[4] &&  s[3] &&          !s[1] &&  s[0] &&  d[3] &&  d[2] &&  d[1])            ||
// 				( !s[4] &&  s[3] &&          !s[1] &&  s[0] &&  d[3] &&  d[2] &&           d[0])   ||
// 				( !s[4] &&  s[3] &&          !s[1] && !s[0] &&  d[3] &&  d[2] && !d[1])            ||
// 				( !s[4] &&  s[3] &&                    s[0] &&  d[3] &&  d[2] &&  d[1] &&  d[0])   ||
// 				( !s[4] && !s[3] &&  s[2] &&  s[1] &&  s[0] &&  d[3] && !d[2] )                    ||
// 				( !s[4] && !s[3] &&  s[2] &&  s[1] &&  s[0] &&  d[3] &&          !d[1] && !d[0])   ||
// 				( !s[4] && !s[3] &&  s[2] &&  s[1] &&           d[3] && !d[2] && !d[1])            ||
// 				( !s[4] && !s[3] &&  s[2] &&  s[1] &&           d[3] && !d[2] &&          !d[0]) ;

// updated
assign mul_3 = 
( !s[4]  &&  s[3]  &&  s[2] &&          !s[0] &&  d[3] &&  d[2] &&  d[1])         ||
( !s[4]  &&  s[3]  && !s[2] &&  s[1] &&           d[3] &&  d[2])                  ||
( !s[4]  &&  s[3]  && !s[2] && !s[1] &&           d[3] &&           d[1] && !d[0])||
( !s[4]  &&  s[3]  && !s[2] && !s[1] &&           d[3] &&          !d[1] &&  d[0])||
( !s[4]  &&  s[3]  && !s[2] &&           s[0] &&  d[3] &&  d[2])                  ||
( !s[4]  &&  s[3]  && !s[2] &&          !s[0] &&  d[3] &&          !d[1] && !d[0])||
( !s[4]  &&  s[3]  && !s[2] &&                    d[3] && !d[2] &&  d[1] &&  d[0])||
( !s[4]  &&  s[3]  &&          !s[1] &&  s[0] &&  d[3] &&  d[2] &&  d[1])         ||
( !s[4]  &&  s[3]  &&          !s[1] && !s[0] &&  d[3] &&  d[2] && !d[1])         ||
( !s[4]  &&  s[3]  &&          !s[1] &&           d[3] &&  d[2] && !d[1] &&  d[0])||
( !s[4]  &&  s[3]  &&                    s[0] &&  d[3] &&  d[2] &&  d[1] &&  d[0])||
( !s[4]  && !s[3]  &&  s[2] &&  s[1] &&  s[0] &&  d[3] && !d[2])                  ||
( !s[4]  && !s[3]  &&  s[2] &&  s[1] &&  s[0] &&  d[3] &&          !d[1]&&  !d[0])||
( !s[4]  && !s[3]  &&  s[2] &&  s[1] &&           d[3] && !d[2] && !d[1])         ||
( !s[4]  && !s[3]  &&  s[2] &&  s[1] &&           d[3] && !d[2] &&          !d[0])||
( !s[4]  && !s[3]  &&  s[2] &&           s[0] &&  d[3] && !d[2] && !d[1]) ;


endmodule
