module Division_tb();

	reg [31:0] inA,inB;
	reg clk,en,n_rst;
	wire [31:0] out;
	wire finish;

Division DV(inA,inB,clk,en,n_rst,out,finish);


initial begin
	clk = 0 ;
	en = 1 ;
	n_rst = 0 ;

	//Normal cases
	inA=32'b01000010111010000000000000000000; inB=32'b01000000010000000000000000000000; //116 / 3
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01000010111010000000000000000000; inB=32'b11000000010000000000000000000000; //116 / (-3)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11000010111010000000000000000000; inB=32'b01000000010000000000000000000000; //-116 / 3
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11000010111010000000000000000000; inB=32'b11000000010000000000000000000000; //-116 / (-3)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b01000010111101101110100101111001; //0.69 / 123.456
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b11000010111101101110100101111001; //0.69 / (-123.456)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b01000010111101101110100101111001; //-0.69 / 123.456
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b11000010111101101110100101111001; //-0.69 / (-123.456)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b00111111001100001010001111010111; //0.69 / 0.69
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11000010111010000000000000000000; inB=32'b11000010111010000000000000000000; //-116 / (-116)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;

	//Zero cases
	inA=32'b00000000000000000000000000000000; inB=32'b01000000010000000000000000000000;
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01000000010000000000000000000000; // 0 / 3
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b11000000010000000000000000000000;
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b11000000010000000000000000000000; // 0 / (-3)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b00000000000000000000000000000000;
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b10000000000000000000000000000000; // 0.69 / 0
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b00000000000000000000000000000000;
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b10000000000000000000000000000000; // -0.69 / 0
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b10000000000000000000000000000000;
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b00000000000000000000000000000000;
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b10000000000000000000000000000000; // 0 / 0
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;

	//Infinity cases
	inA=32'b01111111100000000000000000000000; inB=32'b01000000010000000000000000000000;	// inf / 3
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01000000010000000000000000000000; // -inf / 3
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b11000000010000000000000000000000;	// inf / (-3)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b11000000010000000000000000000000; // -inf / (-3)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b01111111100000000000000000000000;	// 0.69 / inf
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b11111111100000000000000000000000; // 0.69 / (-inf)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b01111111100000000000000000000000;	// -0.69 / inf
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b11111111100000000000000000000000; // -0.69 / (-inf)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	// inf / inf
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b11111111100000000000000000000000;	// inf / (-inf)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01111111100000000000000000000000;	// -inf / inf
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b11111111100000000000000000000000; // -inf / (-inf)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;

	//Nan cases
	inA=32'b01111111101010101010101010101010; inB=32'b01000000010000000000000000000000;	// NaN / 3
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b11000000010000000000000000000000;	// NaN / (-3)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00111111001100001010001111010111; inB=32'b01111111101010101010101010101010;	// 0.69 / NaN
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10111111001100001010001111010111; inB=32'b01111111101010101010101010101010;	// -0.69 / NaN
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b01111111101010101010101010101010;	// NaN / NaN
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;

	//Crossover
	inA=32'b00000000000000000000000000000000; inB=32'b01111111100000000000000000000000;	
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01111111100000000000000000000000; // 0 / inf
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b11111111100000000000000000000000;	
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b11111111100000000000000000000000; // 0 / (-inf)
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b00000000000000000000000000000000; inB=32'b01111111101010101010101010101010;	
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b10000000000000000000000000000000; inB=32'b01111111101010101010101010101010; // 0 / NaN
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b00000000000000000000000000000000;	
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b10000000000000000000000000000000; // inf / 0
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b00000000000000000000000000000000;	
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b10000000000000000000000000000000; // -inf / 0
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111100000000000000000000000; inB=32'b01111111101010101010101010101010;	// inf / NaN
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b11111111100000000000000000000000; inB=32'b01111111101010101010101010101010; // -inf / NaN
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b00000000000000000000000000000000;	
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b10000000000000000000000000000000; // NaN / 0
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b01111111100000000000000000000000;	// NaN / inf
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	inA=32'b01111111101010101010101010101010; inB=32'b11111111100000000000000000000000; // NaN / (-inf)m
	#20 n_rst = 1 ; #260 ; n_rst = 0 ;
	$finish ;
end


always begin
	clk=~clk ;
	#10 ;
end


endmodule


